VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CF_SRAM_1024x32
  CLASS BLOCK ;
  FOREIGN CF_SRAM_1024x32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 387.870 BY 306.775 ;
  PIN WLOFF
    PORT
      LAYER met1 ;
        RECT 193.805 306.055 194.065 306.775 ;
        RECT 203.450 3.000 203.705 3.675 ;
        RECT 203.445 0.000 203.705 3.000 ;
      LAYER met2 ;
        RECT 193.750 306.465 194.120 306.745 ;
        RECT 193.750 2.420 194.120 2.490 ;
        RECT 203.415 2.420 203.735 2.480 ;
        RECT 193.750 2.280 203.735 2.420 ;
        RECT 193.750 2.210 194.120 2.280 ;
        RECT 203.415 2.220 203.735 2.280 ;
      LAYER met3 ;
        RECT 193.770 306.440 194.100 306.770 ;
        RECT 193.785 2.515 194.085 306.440 ;
        RECT 193.770 2.185 194.100 2.515 ;
    END
  END WLOFF
  PIN DO[16]
    PORT
      LAYER met1 ;
        RECT 211.405 0.000 211.635 3.500 ;
    END
  END DO[16]
  PIN BEN[16]
    PORT
      LAYER met1 ;
        RECT 217.545 0.000 217.775 3.500 ;
    END
  END BEN[16]
  PIN DO[17]
    PORT
      LAYER met1 ;
        RECT 222.305 0.000 222.535 3.500 ;
    END
  END DO[17]
  PIN BEN[17]
    PORT
      LAYER met1 ;
        RECT 228.445 0.000 228.675 3.500 ;
    END
  END BEN[17]
  PIN DO[18]
    PORT
      LAYER met1 ;
        RECT 233.205 0.000 233.435 3.500 ;
    END
  END DO[18]
  PIN BEN[18]
    PORT
      LAYER met1 ;
        RECT 239.345 0.000 239.575 3.500 ;
    END
  END BEN[18]
  PIN DO[19]
    PORT
      LAYER met1 ;
        RECT 244.105 0.000 244.335 3.500 ;
    END
  END DO[19]
  PIN BEN[19]
    PORT
      LAYER met1 ;
        RECT 250.245 0.000 250.475 3.500 ;
    END
  END BEN[19]
  PIN DO[20]
    PORT
      LAYER met1 ;
        RECT 255.005 0.000 255.235 3.500 ;
    END
  END DO[20]
  PIN BEN[20]
    PORT
      LAYER met1 ;
        RECT 261.145 0.000 261.375 3.500 ;
    END
  END BEN[20]
  PIN DO[21]
    PORT
      LAYER met1 ;
        RECT 265.905 0.000 266.135 3.500 ;
    END
  END DO[21]
  PIN BEN[21]
    PORT
      LAYER met1 ;
        RECT 272.045 0.000 272.275 3.500 ;
    END
  END BEN[21]
  PIN DO[22]
    PORT
      LAYER met1 ;
        RECT 276.805 0.000 277.035 3.500 ;
    END
  END DO[22]
  PIN BEN[22]
    PORT
      LAYER met1 ;
        RECT 282.945 0.000 283.175 3.500 ;
    END
  END BEN[22]
  PIN DO[23]
    PORT
      LAYER met1 ;
        RECT 287.705 0.000 287.935 3.500 ;
    END
  END DO[23]
  PIN BEN[23]
    PORT
      LAYER met1 ;
        RECT 293.845 0.000 294.075 3.500 ;
    END
  END BEN[23]
  PIN DO[24]
    PORT
      LAYER met1 ;
        RECT 298.605 0.000 298.835 3.500 ;
    END
  END DO[24]
  PIN BEN[24]
    PORT
      LAYER met1 ;
        RECT 304.745 0.000 304.975 3.500 ;
    END
  END BEN[24]
  PIN DO[25]
    PORT
      LAYER met1 ;
        RECT 309.505 0.000 309.735 3.500 ;
    END
  END DO[25]
  PIN BEN[25]
    PORT
      LAYER met1 ;
        RECT 315.645 0.000 315.875 3.500 ;
    END
  END BEN[25]
  PIN DO[26]
    PORT
      LAYER met1 ;
        RECT 320.405 0.000 320.635 3.500 ;
    END
  END DO[26]
  PIN BEN[26]
    PORT
      LAYER met1 ;
        RECT 326.545 0.000 326.775 3.500 ;
    END
  END BEN[26]
  PIN DO[27]
    PORT
      LAYER met1 ;
        RECT 331.305 0.000 331.535 3.500 ;
    END
  END DO[27]
  PIN BEN[27]
    PORT
      LAYER met1 ;
        RECT 337.445 0.000 337.675 3.500 ;
    END
  END BEN[27]
  PIN DO[28]
    PORT
      LAYER met1 ;
        RECT 342.205 0.000 342.435 3.500 ;
    END
  END DO[28]
  PIN BEN[28]
    PORT
      LAYER met1 ;
        RECT 348.345 0.000 348.575 3.500 ;
    END
  END BEN[28]
  PIN DO[29]
    PORT
      LAYER met1 ;
        RECT 353.105 0.000 353.335 3.500 ;
    END
  END DO[29]
  PIN BEN[29]
    PORT
      LAYER met1 ;
        RECT 359.245 0.000 359.475 3.500 ;
    END
  END BEN[29]
  PIN DO[30]
    PORT
      LAYER met1 ;
        RECT 364.005 0.000 364.235 3.500 ;
    END
  END DO[30]
  PIN BEN[30]
    PORT
      LAYER met1 ;
        RECT 370.145 0.000 370.375 3.500 ;
    END
  END BEN[30]
  PIN DO[31]
    PORT
      LAYER met1 ;
        RECT 374.905 0.000 375.135 3.500 ;
    END
  END DO[31]
  PIN BEN[31]
    PORT
      LAYER met1 ;
        RECT 381.045 0.000 381.275 3.500 ;
    END
  END BEN[31]
  PIN AD[0]
    PORT
      LAYER met1 ;
        RECT 199.905 0.000 200.165 3.510 ;
    END
  END AD[0]
  PIN AD[1]
    PORT
      LAYER met1 ;
        RECT 196.765 0.000 197.025 3.510 ;
    END
  END AD[1]
  PIN AD[2]
    PORT
      LAYER met1 ;
        RECT 196.365 0.000 196.625 3.510 ;
    END
  END AD[2]
  PIN WLBI
    PORT
      LAYER met1 ;
        RECT 220.735 0.000 220.975 3.635 ;
    END
  END WLBI
  PIN CLKin
    PORT
      LAYER met1 ;
        RECT 227.045 0.000 227.275 3.645 ;
    END
  END CLKin
  PIN EN
    PORT
      LAYER met1 ;
        RECT 203.845 0.000 204.105 3.665 ;
    END
  END EN
  PIN R_WB
    PORT
      LAYER met1 ;
        RECT 200.305 0.000 200.565 3.505 ;
    END
  END R_WB
  PIN SM
    PORT
      LAYER met1 ;
        RECT 208.185 0.000 208.385 3.865 ;
    END
  END SM
  PIN TM
    PORT
      LAYER met1 ;
        RECT 220.345 0.000 220.595 3.630 ;
    END
  END TM
  PIN ScanInDR
    PORT
      LAYER met1 ;
        RECT 209.885 0.000 210.075 3.785 ;
    END
  END ScanInDR
  PIN ScanOutCC
    PORT
      LAYER met1 ;
        RECT 208.525 0.000 208.725 3.880 ;
    END
  END ScanOutCC
  PIN ScanInDL
    PORT
      LAYER met1 ;
        RECT 171.915 0.000 172.105 4.015 ;
    END
  END ScanInDL
  PIN DO[9]
    PORT
      LAYER met1 ;
        RECT 78.135 0.000 78.365 3.500 ;
    END
  END DO[9]
  PIN BEN[9]
    PORT
      LAYER met1 ;
        RECT 71.995 0.000 72.225 3.500 ;
    END
  END BEN[9]
  PIN DO[10]
    PORT
      LAYER met1 ;
        RECT 67.235 0.000 67.465 3.500 ;
    END
  END DO[10]
  PIN BEN[10]
    PORT
      LAYER met1 ;
        RECT 61.095 0.000 61.325 3.500 ;
    END
  END BEN[10]
  PIN DO[11]
    PORT
      LAYER met1 ;
        RECT 56.335 0.000 56.565 3.500 ;
    END
  END DO[11]
  PIN BEN[11]
    PORT
      LAYER met1 ;
        RECT 50.195 0.000 50.425 3.500 ;
    END
  END BEN[11]
  PIN DO[12]
    PORT
      LAYER met1 ;
        RECT 45.435 0.000 45.665 3.500 ;
    END
  END DO[12]
  PIN BEN[12]
    PORT
      LAYER met1 ;
        RECT 39.295 0.000 39.525 3.500 ;
    END
  END BEN[12]
  PIN DO[13]
    PORT
      LAYER met1 ;
        RECT 34.535 0.000 34.765 3.500 ;
    END
  END DO[13]
  PIN BEN[13]
    PORT
      LAYER met1 ;
        RECT 28.395 0.000 28.625 3.500 ;
    END
  END BEN[13]
  PIN DO[14]
    PORT
      LAYER met1 ;
        RECT 23.635 0.000 23.865 3.500 ;
    END
  END DO[14]
  PIN BEN[14]
    PORT
      LAYER met1 ;
        RECT 17.495 0.000 17.725 3.500 ;
    END
  END BEN[14]
  PIN DO[15]
    PORT
      LAYER met1 ;
        RECT 12.735 0.000 12.965 3.500 ;
    END
  END DO[15]
  PIN BEN[15]
    PORT
      LAYER met1 ;
        RECT 6.595 0.000 6.825 3.500 ;
    END
  END BEN[15]
  PIN BEN[8]
    PORT
      LAYER met1 ;
        RECT 82.895 0.000 83.125 3.500 ;
    END
  END BEN[8]
  PIN AD[3]
    PORT
      LAYER met1 ;
        RECT 179.065 0.000 179.325 3.620 ;
    END
  END AD[3]
  PIN AD[4]
    PORT
      LAYER met1 ;
        RECT 189.685 0.000 189.945 3.575 ;
    END
  END AD[4]
  PIN AD[5]
    PORT
      LAYER met1 ;
        RECT 189.285 0.000 189.545 3.000 ;
    END
  END AD[5]
  PIN AD[6]
    PORT
      LAYER met1 ;
        RECT 186.145 0.000 186.405 3.535 ;
    END
  END AD[6]
  PIN AD[7]
    PORT
      LAYER met1 ;
        RECT 185.745 0.000 186.005 3.000 ;
    END
  END AD[7]
  PIN AD[8]
    PORT
      LAYER met1 ;
        RECT 182.605 0.000 182.865 3.610 ;
    END
  END AD[8]
  PIN AD[9]
    PORT
      LAYER met1 ;
        RECT 182.205 0.000 182.465 3.605 ;
    END
  END AD[9]
  PIN ScanInCC
    PORT
      LAYER met1 ;
        RECT 178.140 0.000 178.400 3.630 ;
    END
  END ScanInCC
  PIN DO[0]
    PORT
      LAYER met1 ;
        RECT 176.235 0.000 176.465 3.500 ;
    END
  END DO[0]
  PIN BEN[0]
    PORT
      LAYER met1 ;
        RECT 170.095 0.000 170.325 3.500 ;
    END
  END BEN[0]
  PIN DO[1]
    PORT
      LAYER met1 ;
        RECT 165.335 0.000 165.565 3.500 ;
    END
  END DO[1]
  PIN BEN[1]
    PORT
      LAYER met1 ;
        RECT 159.195 0.000 159.425 3.500 ;
    END
  END BEN[1]
  PIN DO[2]
    PORT
      LAYER met1 ;
        RECT 154.435 0.000 154.665 3.500 ;
    END
  END DO[2]
  PIN BEN[2]
    PORT
      LAYER met1 ;
        RECT 148.295 0.000 148.525 3.500 ;
    END
  END BEN[2]
  PIN DO[3]
    PORT
      LAYER met1 ;
        RECT 143.535 0.000 143.765 3.500 ;
    END
  END DO[3]
  PIN BEN[3]
    PORT
      LAYER met1 ;
        RECT 137.395 0.000 137.625 3.500 ;
    END
  END BEN[3]
  PIN DO[4]
    PORT
      LAYER met1 ;
        RECT 132.635 0.000 132.865 3.500 ;
    END
  END DO[4]
  PIN BEN[4]
    PORT
      LAYER met1 ;
        RECT 126.495 0.000 126.725 3.500 ;
    END
  END BEN[4]
  PIN DO[5]
    PORT
      LAYER met1 ;
        RECT 121.735 0.000 121.965 3.500 ;
    END
  END DO[5]
  PIN BEN[5]
    PORT
      LAYER met1 ;
        RECT 115.595 0.000 115.825 3.500 ;
    END
  END BEN[5]
  PIN DO[6]
    PORT
      LAYER met1 ;
        RECT 110.835 0.000 111.065 3.500 ;
    END
  END DO[6]
  PIN BEN[6]
    PORT
      LAYER met1 ;
        RECT 104.695 0.000 104.925 3.500 ;
    END
  END BEN[6]
  PIN DO[7]
    PORT
      LAYER met1 ;
        RECT 99.935 0.000 100.165 3.500 ;
    END
  END DO[7]
  PIN BEN[7]
    PORT
      LAYER met1 ;
        RECT 93.795 0.000 94.025 3.500 ;
    END
  END BEN[7]
  PIN DO[8]
    PORT
      LAYER met1 ;
        RECT 89.035 0.000 89.265 3.500 ;
    END
  END DO[8]
  PIN DI[3]
    PORT
      LAYER met1 ;
        RECT 142.275 0.000 142.505 3.430 ;
    END
  END DI[3]
  PIN DI[12]
    PORT
      LAYER met1 ;
        RECT 44.175 0.000 44.405 3.430 ;
    END
  END DI[12]
  PIN DI[0]
    PORT
      LAYER met1 ;
        RECT 174.975 0.000 175.205 3.430 ;
    END
  END DI[0]
  PIN DI[4]
    PORT
      LAYER met1 ;
        RECT 131.375 0.000 131.605 3.430 ;
    END
  END DI[4]
  PIN DI[14]
    PORT
      LAYER met1 ;
        RECT 22.375 0.000 22.605 3.430 ;
    END
  END DI[14]
  PIN DI[11]
    PORT
      LAYER met1 ;
        RECT 55.075 0.000 55.305 3.430 ;
    END
  END DI[11]
  PIN DI[5]
    PORT
      LAYER met1 ;
        RECT 120.475 0.000 120.705 3.430 ;
    END
  END DI[5]
  PIN DI[1]
    PORT
      LAYER met1 ;
        RECT 164.075 0.000 164.305 3.430 ;
    END
  END DI[1]
  PIN DI[9]
    PORT
      LAYER met1 ;
        RECT 76.875 0.000 77.105 3.430 ;
    END
  END DI[9]
  PIN DI[6]
    PORT
      LAYER met1 ;
        RECT 109.575 0.000 109.805 3.430 ;
    END
  END DI[6]
  PIN DI[15]
    PORT
      LAYER met1 ;
        RECT 11.475 0.000 11.705 3.430 ;
    END
  END DI[15]
  PIN DI[2]
    PORT
      LAYER met1 ;
        RECT 153.175 0.000 153.405 3.430 ;
    END
  END DI[2]
  PIN DI[7]
    PORT
      LAYER met1 ;
        RECT 98.675 0.000 98.905 3.430 ;
    END
  END DI[7]
  PIN DI[13]
    PORT
      LAYER met1 ;
        RECT 33.275 0.000 33.505 3.430 ;
    END
  END DI[13]
  PIN DI[10]
    PORT
      LAYER met1 ;
        RECT 65.975 0.000 66.205 3.430 ;
    END
  END DI[10]
  PIN DI[8]
    PORT
      LAYER met1 ;
        RECT 87.775 0.000 88.005 3.430 ;
    END
  END DI[8]
  PIN DI[23]
    PORT
      LAYER met1 ;
        RECT 288.965 0.000 289.195 3.430 ;
    END
  END DI[23]
  PIN DI[27]
    PORT
      LAYER met1 ;
        RECT 332.565 0.000 332.795 3.430 ;
    END
  END DI[27]
  PIN DI[19]
    PORT
      LAYER met1 ;
        RECT 245.365 0.000 245.595 3.430 ;
    END
  END DI[19]
  PIN DI[21]
    PORT
      LAYER met1 ;
        RECT 267.165 0.000 267.395 3.430 ;
    END
  END DI[21]
  PIN DI[28]
    PORT
      LAYER met1 ;
        RECT 343.465 0.000 343.695 3.430 ;
    END
  END DI[28]
  PIN DI[24]
    PORT
      LAYER met1 ;
        RECT 299.865 0.000 300.095 3.430 ;
    END
  END DI[24]
  PIN DI[18]
    PORT
      LAYER met1 ;
        RECT 234.465 0.000 234.695 3.430 ;
    END
  END DI[18]
  PIN DI[29]
    PORT
      LAYER met1 ;
        RECT 354.365 0.000 354.595 3.430 ;
    END
  END DI[29]
  PIN DI[16]
    PORT
      LAYER met1 ;
        RECT 212.665 0.000 212.895 3.430 ;
    END
  END DI[16]
  PIN DI[25]
    PORT
      LAYER met1 ;
        RECT 310.765 0.000 310.995 3.430 ;
    END
  END DI[25]
  PIN DI[30]
    PORT
      LAYER met1 ;
        RECT 365.265 0.000 365.495 3.430 ;
    END
  END DI[30]
  PIN DI[22]
    PORT
      LAYER met1 ;
        RECT 278.065 0.000 278.295 3.430 ;
    END
  END DI[22]
  PIN DI[20]
    PORT
      LAYER met1 ;
        RECT 256.265 0.000 256.495 3.430 ;
    END
  END DI[20]
  PIN DI[26]
    PORT
      LAYER met1 ;
        RECT 321.665 0.000 321.895 3.430 ;
    END
  END DI[26]
  PIN DI[17]
    PORT
      LAYER met1 ;
        RECT 223.565 0.000 223.795 3.430 ;
    END
  END DI[17]
  PIN DI[31]
    PORT
      LAYER met1 ;
        RECT 376.165 0.000 376.395 3.430 ;
    END
  END DI[31]
  PIN vnb
    PORT
      LAYER met2 ;
        RECT 1.230 273.890 386.640 274.360 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 259.440 386.640 259.910 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 244.990 386.640 245.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 230.540 386.640 231.010 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 216.090 386.640 216.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 201.640 386.640 202.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 187.190 386.640 187.660 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 172.740 386.640 173.210 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 158.290 386.640 158.760 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 288.340 386.640 288.810 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 143.840 386.640 144.310 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 129.390 386.640 129.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 114.940 386.640 115.410 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 100.490 386.640 100.960 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.230 86.040 386.640 86.510 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 46.925 178.430 47.565 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 14.355 383.840 14.935 ;
        RECT 4.030 14.295 178.430 14.355 ;
        RECT 209.440 14.295 383.840 14.355 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 13.355 0.960 14.935 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 13.355 387.870 14.935 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.440 46.925 383.840 47.565 ;
    END
  END vnb
  PIN vpwrm
    PORT
      LAYER met2 ;
        RECT 4.030 15.865 383.840 16.745 ;
        RECT 4.030 15.745 178.430 15.865 ;
        RECT 209.440 15.745 383.840 15.865 ;
    END
  END vpwrm
  PIN vpwra
    PORT
      LAYER met2 ;
        RECT 1.780 304.655 386.090 305.655 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.780 72.040 179.080 72.510 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 52.260 0.960 54.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 19.895 383.840 20.595 ;
    END
    PORT
      LAYER met2 ;
        RECT 208.790 72.040 386.090 72.510 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 52.260 387.870 54.440 ;
    END
  END vpwra
  PIN vpwrp
    PORT
      LAYER met2 ;
        RECT 0.980 67.265 179.080 68.265 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 57.860 0.980 66.205 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 51.175 178.430 51.815 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 48.605 383.840 49.245 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 42.015 383.840 42.655 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 39.535 0.960 41.645 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 39.050 383.840 39.690 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 33.320 383.840 33.960 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 25.810 383.840 26.710 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 24.310 0.960 25.890 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 19.165 383.840 19.745 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 16.895 383.840 17.475 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 4.010 383.840 4.880 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 3.360 0.960 4.935 ;
    END
    PORT
      LAYER met2 ;
        RECT 208.790 67.265 386.890 68.265 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 24.310 387.870 25.890 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.890 57.860 387.870 66.205 ;
    END
    PORT
      LAYER met2 ;
        RECT 209.440 51.175 383.840 51.815 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 3.360 387.870 4.935 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 39.535 387.870 41.645 ;
    END
  END vpwrp
  PIN vgnd
    PORT
      LAYER met2 ;
        RECT 387.590 304.050 387.870 306.315 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.140 305.795 386.730 306.315 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 304.050 0.280 306.315 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.140 71.000 179.080 71.470 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 54.815 383.840 55.365 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 47.765 383.840 48.405 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 45.065 0.960 48.840 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 43.205 383.840 43.845 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 41.285 383.840 41.865 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 37.675 383.840 38.315 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 34.785 383.840 35.425 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 32.590 383.840 33.170 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 31.070 383.840 31.650 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 29.310 0.960 30.890 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 26.860 383.840 27.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 178.430 24.370 209.440 24.690 ;
        RECT 4.030 24.110 383.840 24.370 ;
        RECT 4.030 23.790 178.430 24.110 ;
        RECT 209.440 23.790 383.840 24.110 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 20.745 383.840 21.325 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 13.565 383.840 14.145 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 8.355 0.960 9.935 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 3.000 383.840 3.870 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 45.065 387.870 48.840 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 29.310 387.870 30.890 ;
    END
    PORT
      LAYER met2 ;
        RECT 208.790 71.000 386.730 71.470 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 8.355 387.870 9.935 ;
    END
  END vgnd
  PIN vpb
    PORT
      LAYER met2 ;
        RECT 3.010 289.075 384.860 289.545 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 274.625 384.860 275.095 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 260.175 384.860 260.645 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 245.725 384.860 246.195 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 231.275 384.860 231.745 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 216.825 384.860 217.295 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 202.375 384.860 202.845 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 187.925 384.860 188.395 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 173.475 384.860 173.945 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 159.025 384.860 159.495 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 144.575 384.860 145.045 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 130.125 384.860 130.595 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 115.675 384.860 116.145 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 101.225 384.860 101.695 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.010 86.775 384.860 87.245 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.900 50.385 383.970 51.025 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.000 34.310 0.960 36.115 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.030 17.625 383.840 18.205 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 34.310 387.870 36.115 ;
    END
  END vpb
  PIN vpwrpc
    PORT
      LAYER met2 ;
        RECT 0.000 18.355 0.960 18.615 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 18.355 387.870 18.615 ;
    END
  END vpwrpc
  PIN vpwrac
    PORT
      LAYER met2 ;
        RECT 0.000 20.235 0.960 20.495 ;
    END
    PORT
      LAYER met2 ;
        RECT 386.910 20.235 387.870 20.495 ;
    END
  END vpwrac
  OBS
      LAYER li1 ;
        RECT 0.000 3.000 387.870 306.315 ;
      LAYER met1 ;
        RECT 0.000 306.035 1.140 306.315 ;
      LAYER met1 ;
        RECT 1.140 306.035 2.835 306.315 ;
      LAYER met1 ;
        RECT 2.835 306.035 5.080 306.315 ;
        RECT 0.000 305.980 5.080 306.035 ;
      LAYER met1 ;
        RECT 5.080 305.980 5.580 306.315 ;
      LAYER met1 ;
        RECT 5.580 306.035 13.370 306.315 ;
      LAYER met1 ;
        RECT 13.370 306.035 15.610 306.315 ;
      LAYER met1 ;
        RECT 15.610 306.055 193.805 306.315 ;
        RECT 194.065 306.055 372.260 306.315 ;
        RECT 15.610 306.035 372.260 306.055 ;
      LAYER met1 ;
        RECT 372.260 306.035 374.500 306.315 ;
      LAYER met1 ;
        RECT 374.500 306.035 382.290 306.315 ;
        RECT 5.580 305.980 382.290 306.035 ;
      LAYER met1 ;
        RECT 382.290 305.980 382.790 306.315 ;
      LAYER met1 ;
        RECT 382.790 306.035 385.035 306.315 ;
      LAYER met1 ;
        RECT 385.035 306.035 386.730 306.315 ;
      LAYER met1 ;
        RECT 386.730 306.035 387.870 306.315 ;
        RECT 382.790 305.980 387.870 306.035 ;
        RECT 0.000 4.015 387.870 305.980 ;
        RECT 0.000 4.000 171.915 4.015 ;
        RECT 0.000 3.500 8.745 4.000 ;
        RECT 0.000 3.000 6.595 3.500 ;
        RECT 6.825 3.000 8.745 3.500 ;
      LAYER met1 ;
        RECT 8.745 3.000 10.115 4.000 ;
      LAYER met1 ;
        RECT 10.115 3.500 19.645 4.000 ;
        RECT 10.115 3.430 12.735 3.500 ;
        RECT 10.115 3.000 11.475 3.430 ;
        RECT 11.705 3.000 12.735 3.430 ;
        RECT 12.965 3.000 17.495 3.500 ;
        RECT 17.725 3.000 19.645 3.500 ;
      LAYER met1 ;
        RECT 19.645 3.000 21.015 4.000 ;
      LAYER met1 ;
        RECT 21.015 3.500 30.545 4.000 ;
        RECT 21.015 3.430 23.635 3.500 ;
        RECT 21.015 3.000 22.375 3.430 ;
        RECT 22.605 3.000 23.635 3.430 ;
        RECT 23.865 3.000 28.395 3.500 ;
        RECT 28.625 3.000 30.545 3.500 ;
      LAYER met1 ;
        RECT 30.545 3.000 31.915 4.000 ;
      LAYER met1 ;
        RECT 31.915 3.500 41.445 4.000 ;
        RECT 31.915 3.430 34.535 3.500 ;
        RECT 31.915 3.000 33.275 3.430 ;
        RECT 33.505 3.000 34.535 3.430 ;
        RECT 34.765 3.000 39.295 3.500 ;
        RECT 39.525 3.000 41.445 3.500 ;
      LAYER met1 ;
        RECT 41.445 3.000 42.815 4.000 ;
      LAYER met1 ;
        RECT 42.815 3.500 52.345 4.000 ;
        RECT 42.815 3.430 45.435 3.500 ;
        RECT 42.815 3.000 44.175 3.430 ;
        RECT 44.405 3.000 45.435 3.430 ;
        RECT 45.665 3.000 50.195 3.500 ;
        RECT 50.425 3.000 52.345 3.500 ;
      LAYER met1 ;
        RECT 52.345 3.000 53.715 4.000 ;
      LAYER met1 ;
        RECT 53.715 3.500 63.245 4.000 ;
        RECT 53.715 3.430 56.335 3.500 ;
        RECT 53.715 3.000 55.075 3.430 ;
        RECT 55.305 3.000 56.335 3.430 ;
        RECT 56.565 3.000 61.095 3.500 ;
        RECT 61.325 3.000 63.245 3.500 ;
      LAYER met1 ;
        RECT 63.245 3.000 64.615 4.000 ;
      LAYER met1 ;
        RECT 64.615 3.500 74.145 4.000 ;
        RECT 64.615 3.430 67.235 3.500 ;
        RECT 64.615 3.000 65.975 3.430 ;
        RECT 66.205 3.000 67.235 3.430 ;
        RECT 67.465 3.000 71.995 3.500 ;
        RECT 72.225 3.000 74.145 3.500 ;
      LAYER met1 ;
        RECT 74.145 3.000 75.515 4.000 ;
      LAYER met1 ;
        RECT 75.515 3.500 85.045 4.000 ;
        RECT 75.515 3.430 78.135 3.500 ;
        RECT 75.515 3.000 76.875 3.430 ;
        RECT 77.105 3.000 78.135 3.430 ;
        RECT 78.365 3.000 82.895 3.500 ;
        RECT 83.125 3.000 85.045 3.500 ;
      LAYER met1 ;
        RECT 85.045 3.000 86.415 4.000 ;
      LAYER met1 ;
        RECT 86.415 3.500 95.945 4.000 ;
        RECT 86.415 3.430 89.035 3.500 ;
        RECT 86.415 3.000 87.775 3.430 ;
        RECT 88.005 3.000 89.035 3.430 ;
        RECT 89.265 3.000 93.795 3.500 ;
        RECT 94.025 3.000 95.945 3.500 ;
      LAYER met1 ;
        RECT 95.945 3.000 97.315 4.000 ;
      LAYER met1 ;
        RECT 97.315 3.500 106.845 4.000 ;
        RECT 97.315 3.430 99.935 3.500 ;
        RECT 97.315 3.000 98.675 3.430 ;
        RECT 98.905 3.000 99.935 3.430 ;
        RECT 100.165 3.000 104.695 3.500 ;
        RECT 104.925 3.000 106.845 3.500 ;
      LAYER met1 ;
        RECT 106.845 3.000 108.215 4.000 ;
      LAYER met1 ;
        RECT 108.215 3.500 117.745 4.000 ;
        RECT 108.215 3.430 110.835 3.500 ;
        RECT 108.215 3.000 109.575 3.430 ;
        RECT 109.805 3.000 110.835 3.430 ;
        RECT 111.065 3.000 115.595 3.500 ;
        RECT 115.825 3.000 117.745 3.500 ;
      LAYER met1 ;
        RECT 117.745 3.000 119.115 4.000 ;
      LAYER met1 ;
        RECT 119.115 3.500 128.645 4.000 ;
        RECT 119.115 3.430 121.735 3.500 ;
        RECT 119.115 3.000 120.475 3.430 ;
        RECT 120.705 3.000 121.735 3.430 ;
        RECT 121.965 3.000 126.495 3.500 ;
        RECT 126.725 3.000 128.645 3.500 ;
      LAYER met1 ;
        RECT 128.645 3.000 130.015 4.000 ;
      LAYER met1 ;
        RECT 130.015 3.500 139.545 4.000 ;
        RECT 130.015 3.430 132.635 3.500 ;
        RECT 130.015 3.000 131.375 3.430 ;
        RECT 131.605 3.000 132.635 3.430 ;
        RECT 132.865 3.000 137.395 3.500 ;
        RECT 137.625 3.000 139.545 3.500 ;
      LAYER met1 ;
        RECT 139.545 3.000 140.915 4.000 ;
      LAYER met1 ;
        RECT 140.915 3.500 150.445 4.000 ;
        RECT 140.915 3.430 143.535 3.500 ;
        RECT 140.915 3.000 142.275 3.430 ;
        RECT 142.505 3.000 143.535 3.430 ;
        RECT 143.765 3.000 148.295 3.500 ;
        RECT 148.525 3.000 150.445 3.500 ;
      LAYER met1 ;
        RECT 150.445 3.000 151.815 4.000 ;
      LAYER met1 ;
        RECT 151.815 3.500 161.345 4.000 ;
        RECT 151.815 3.430 154.435 3.500 ;
        RECT 151.815 3.000 153.175 3.430 ;
        RECT 153.405 3.000 154.435 3.430 ;
        RECT 154.665 3.000 159.195 3.500 ;
        RECT 159.425 3.000 161.345 3.500 ;
      LAYER met1 ;
        RECT 161.345 3.000 162.715 4.000 ;
      LAYER met1 ;
        RECT 162.715 3.500 171.915 4.000 ;
        RECT 162.715 3.430 165.335 3.500 ;
        RECT 162.715 3.000 164.075 3.430 ;
        RECT 164.305 3.000 165.335 3.430 ;
        RECT 165.565 3.000 170.095 3.500 ;
        RECT 170.325 3.000 171.915 3.500 ;
        RECT 172.105 4.000 387.870 4.015 ;
        RECT 172.105 3.000 172.245 4.000 ;
      LAYER met1 ;
        RECT 172.245 3.000 173.615 4.000 ;
      LAYER met1 ;
        RECT 173.615 3.880 214.255 4.000 ;
        RECT 173.615 3.865 208.525 3.880 ;
        RECT 173.615 3.675 208.185 3.865 ;
        RECT 173.615 3.630 203.450 3.675 ;
        RECT 173.615 3.500 178.140 3.630 ;
        RECT 173.615 3.430 176.235 3.500 ;
        RECT 173.615 3.000 174.975 3.430 ;
        RECT 175.205 3.000 176.235 3.430 ;
        RECT 176.465 3.000 178.140 3.500 ;
        RECT 178.400 3.620 203.450 3.630 ;
        RECT 178.400 3.000 179.065 3.620 ;
        RECT 179.325 3.610 203.450 3.620 ;
        RECT 179.325 3.605 182.605 3.610 ;
        RECT 179.325 3.000 182.205 3.605 ;
        RECT 182.465 3.000 182.605 3.605 ;
        RECT 182.865 3.590 203.450 3.610 ;
        RECT 182.865 3.550 189.285 3.590 ;
        RECT 182.865 3.005 185.745 3.550 ;
      LAYER met1 ;
        RECT 185.745 3.005 186.005 3.550 ;
      LAYER met1 ;
        RECT 186.005 3.535 189.285 3.550 ;
        RECT 186.005 3.005 186.145 3.535 ;
        RECT 182.865 3.000 186.145 3.005 ;
        RECT 186.405 3.005 189.285 3.535 ;
      LAYER met1 ;
        RECT 189.285 3.005 189.545 3.590 ;
      LAYER met1 ;
        RECT 189.545 3.575 203.450 3.590 ;
        RECT 189.545 3.005 189.685 3.575 ;
        RECT 186.405 3.000 189.685 3.005 ;
        RECT 189.945 3.510 203.450 3.575 ;
        RECT 189.945 3.000 196.365 3.510 ;
        RECT 196.625 3.000 196.765 3.510 ;
        RECT 197.025 3.000 199.905 3.510 ;
        RECT 200.165 3.505 203.450 3.510 ;
        RECT 200.165 3.000 200.305 3.505 ;
        RECT 200.565 3.000 203.450 3.505 ;
        RECT 203.705 3.665 208.185 3.675 ;
        RECT 203.705 3.000 203.845 3.665 ;
        RECT 204.105 3.000 208.185 3.665 ;
        RECT 208.385 3.000 208.525 3.865 ;
        RECT 208.725 3.785 214.255 3.880 ;
        RECT 208.725 3.000 209.885 3.785 ;
        RECT 210.075 3.500 214.255 3.785 ;
        RECT 210.075 3.000 211.405 3.500 ;
        RECT 211.635 3.430 214.255 3.500 ;
        RECT 211.635 3.000 212.665 3.430 ;
        RECT 212.895 3.000 214.255 3.430 ;
      LAYER met1 ;
        RECT 214.255 3.000 215.625 4.000 ;
      LAYER met1 ;
        RECT 215.625 3.635 225.155 4.000 ;
        RECT 215.625 3.630 220.735 3.635 ;
        RECT 215.625 3.500 220.345 3.630 ;
        RECT 215.625 3.000 217.545 3.500 ;
        RECT 217.775 3.000 220.345 3.500 ;
        RECT 220.595 3.000 220.735 3.630 ;
        RECT 220.975 3.500 225.155 3.635 ;
        RECT 220.975 3.000 222.305 3.500 ;
        RECT 222.535 3.430 225.155 3.500 ;
        RECT 222.535 3.000 223.565 3.430 ;
        RECT 223.795 3.000 225.155 3.430 ;
      LAYER met1 ;
        RECT 225.155 3.000 226.525 4.000 ;
      LAYER met1 ;
        RECT 226.525 3.645 236.055 4.000 ;
        RECT 226.525 3.000 227.045 3.645 ;
        RECT 227.275 3.500 236.055 3.645 ;
        RECT 227.275 3.000 228.445 3.500 ;
        RECT 228.675 3.000 233.205 3.500 ;
        RECT 233.435 3.430 236.055 3.500 ;
        RECT 233.435 3.000 234.465 3.430 ;
        RECT 234.695 3.000 236.055 3.430 ;
      LAYER met1 ;
        RECT 236.055 3.000 237.425 4.000 ;
      LAYER met1 ;
        RECT 237.425 3.500 246.955 4.000 ;
        RECT 237.425 3.000 239.345 3.500 ;
        RECT 239.575 3.000 244.105 3.500 ;
        RECT 244.335 3.430 246.955 3.500 ;
        RECT 244.335 3.000 245.365 3.430 ;
        RECT 245.595 3.000 246.955 3.430 ;
      LAYER met1 ;
        RECT 246.955 3.000 248.325 4.000 ;
      LAYER met1 ;
        RECT 248.325 3.500 257.855 4.000 ;
        RECT 248.325 3.000 250.245 3.500 ;
        RECT 250.475 3.000 255.005 3.500 ;
        RECT 255.235 3.430 257.855 3.500 ;
        RECT 255.235 3.000 256.265 3.430 ;
        RECT 256.495 3.000 257.855 3.430 ;
      LAYER met1 ;
        RECT 257.855 3.000 259.225 4.000 ;
      LAYER met1 ;
        RECT 259.225 3.500 268.755 4.000 ;
        RECT 259.225 3.000 261.145 3.500 ;
        RECT 261.375 3.000 265.905 3.500 ;
        RECT 266.135 3.430 268.755 3.500 ;
        RECT 266.135 3.000 267.165 3.430 ;
        RECT 267.395 3.000 268.755 3.430 ;
      LAYER met1 ;
        RECT 268.755 3.000 270.125 4.000 ;
      LAYER met1 ;
        RECT 270.125 3.500 279.655 4.000 ;
        RECT 270.125 3.000 272.045 3.500 ;
        RECT 272.275 3.000 276.805 3.500 ;
        RECT 277.035 3.430 279.655 3.500 ;
        RECT 277.035 3.000 278.065 3.430 ;
        RECT 278.295 3.000 279.655 3.430 ;
      LAYER met1 ;
        RECT 279.655 3.000 281.025 4.000 ;
      LAYER met1 ;
        RECT 281.025 3.500 290.555 4.000 ;
        RECT 281.025 3.000 282.945 3.500 ;
        RECT 283.175 3.000 287.705 3.500 ;
        RECT 287.935 3.430 290.555 3.500 ;
        RECT 287.935 3.000 288.965 3.430 ;
        RECT 289.195 3.000 290.555 3.430 ;
      LAYER met1 ;
        RECT 290.555 3.000 291.925 4.000 ;
      LAYER met1 ;
        RECT 291.925 3.500 301.455 4.000 ;
        RECT 291.925 3.000 293.845 3.500 ;
        RECT 294.075 3.000 298.605 3.500 ;
        RECT 298.835 3.430 301.455 3.500 ;
        RECT 298.835 3.000 299.865 3.430 ;
        RECT 300.095 3.000 301.455 3.430 ;
      LAYER met1 ;
        RECT 301.455 3.000 302.825 4.000 ;
      LAYER met1 ;
        RECT 302.825 3.500 312.355 4.000 ;
        RECT 302.825 3.000 304.745 3.500 ;
        RECT 304.975 3.000 309.505 3.500 ;
        RECT 309.735 3.430 312.355 3.500 ;
        RECT 309.735 3.000 310.765 3.430 ;
        RECT 310.995 3.000 312.355 3.430 ;
      LAYER met1 ;
        RECT 312.355 3.000 313.725 4.000 ;
      LAYER met1 ;
        RECT 313.725 3.500 323.255 4.000 ;
        RECT 313.725 3.000 315.645 3.500 ;
        RECT 315.875 3.000 320.405 3.500 ;
        RECT 320.635 3.430 323.255 3.500 ;
        RECT 320.635 3.000 321.665 3.430 ;
        RECT 321.895 3.000 323.255 3.430 ;
      LAYER met1 ;
        RECT 323.255 3.000 324.625 4.000 ;
      LAYER met1 ;
        RECT 324.625 3.500 334.155 4.000 ;
        RECT 324.625 3.000 326.545 3.500 ;
        RECT 326.775 3.000 331.305 3.500 ;
        RECT 331.535 3.430 334.155 3.500 ;
        RECT 331.535 3.000 332.565 3.430 ;
        RECT 332.795 3.000 334.155 3.430 ;
      LAYER met1 ;
        RECT 334.155 3.000 335.525 4.000 ;
      LAYER met1 ;
        RECT 335.525 3.500 345.055 4.000 ;
        RECT 335.525 3.000 337.445 3.500 ;
        RECT 337.675 3.000 342.205 3.500 ;
        RECT 342.435 3.430 345.055 3.500 ;
        RECT 342.435 3.000 343.465 3.430 ;
        RECT 343.695 3.000 345.055 3.430 ;
      LAYER met1 ;
        RECT 345.055 3.000 346.425 4.000 ;
      LAYER met1 ;
        RECT 346.425 3.500 355.955 4.000 ;
        RECT 346.425 3.000 348.345 3.500 ;
        RECT 348.575 3.000 353.105 3.500 ;
        RECT 353.335 3.430 355.955 3.500 ;
        RECT 353.335 3.000 354.365 3.430 ;
        RECT 354.595 3.000 355.955 3.430 ;
      LAYER met1 ;
        RECT 355.955 3.000 357.325 4.000 ;
      LAYER met1 ;
        RECT 357.325 3.500 366.855 4.000 ;
        RECT 357.325 3.000 359.245 3.500 ;
        RECT 359.475 3.000 364.005 3.500 ;
        RECT 364.235 3.430 366.855 3.500 ;
        RECT 364.235 3.000 365.265 3.430 ;
        RECT 365.495 3.000 366.855 3.430 ;
      LAYER met1 ;
        RECT 366.855 3.000 368.225 4.000 ;
      LAYER met1 ;
        RECT 368.225 3.500 377.755 4.000 ;
        RECT 368.225 3.000 370.145 3.500 ;
        RECT 370.375 3.000 374.905 3.500 ;
        RECT 375.135 3.430 377.755 3.500 ;
        RECT 375.135 3.000 376.165 3.430 ;
        RECT 376.395 3.000 377.755 3.430 ;
      LAYER met1 ;
        RECT 377.755 3.000 379.125 4.000 ;
      LAYER met1 ;
        RECT 379.125 3.500 387.870 4.000 ;
        RECT 379.125 3.000 381.045 3.500 ;
        RECT 381.275 3.000 387.870 3.500 ;
      LAYER met2 ;
        RECT 0.280 305.795 1.140 306.315 ;
        RECT 386.730 305.795 387.590 306.315 ;
        RECT 0.280 305.655 387.590 305.795 ;
        RECT 0.280 304.655 1.780 305.655 ;
        RECT 386.090 304.655 387.590 305.655 ;
        RECT 0.280 304.050 387.590 304.655 ;
        RECT 0.000 289.545 387.870 304.050 ;
        RECT 0.000 289.075 3.010 289.545 ;
        RECT 384.860 289.075 387.870 289.545 ;
        RECT 0.000 288.810 387.870 289.075 ;
        RECT 0.000 288.340 1.230 288.810 ;
        RECT 386.640 288.340 387.870 288.810 ;
        RECT 0.000 275.095 387.870 288.340 ;
        RECT 0.000 274.625 3.010 275.095 ;
        RECT 384.860 274.625 387.870 275.095 ;
        RECT 0.000 274.360 387.870 274.625 ;
        RECT 0.000 273.890 1.230 274.360 ;
        RECT 386.640 273.890 387.870 274.360 ;
        RECT 0.000 260.645 387.870 273.890 ;
        RECT 0.000 260.175 3.010 260.645 ;
        RECT 384.860 260.175 387.870 260.645 ;
        RECT 0.000 259.910 387.870 260.175 ;
        RECT 0.000 259.440 1.230 259.910 ;
        RECT 386.640 259.440 387.870 259.910 ;
        RECT 0.000 246.195 387.870 259.440 ;
        RECT 0.000 245.725 3.010 246.195 ;
        RECT 384.860 245.725 387.870 246.195 ;
        RECT 0.000 245.460 387.870 245.725 ;
        RECT 0.000 244.990 1.230 245.460 ;
        RECT 386.640 244.990 387.870 245.460 ;
        RECT 0.000 231.745 387.870 244.990 ;
        RECT 0.000 231.275 3.010 231.745 ;
        RECT 384.860 231.275 387.870 231.745 ;
        RECT 0.000 231.010 387.870 231.275 ;
        RECT 0.000 230.540 1.230 231.010 ;
        RECT 386.640 230.540 387.870 231.010 ;
        RECT 0.000 217.295 387.870 230.540 ;
        RECT 0.000 216.825 3.010 217.295 ;
        RECT 384.860 216.825 387.870 217.295 ;
        RECT 0.000 216.560 387.870 216.825 ;
        RECT 0.000 216.090 1.230 216.560 ;
        RECT 386.640 216.090 387.870 216.560 ;
        RECT 0.000 202.845 387.870 216.090 ;
        RECT 0.000 202.375 3.010 202.845 ;
        RECT 384.860 202.375 387.870 202.845 ;
        RECT 0.000 202.110 387.870 202.375 ;
        RECT 0.000 201.640 1.230 202.110 ;
        RECT 386.640 201.640 387.870 202.110 ;
        RECT 0.000 188.395 387.870 201.640 ;
        RECT 0.000 187.925 3.010 188.395 ;
        RECT 384.860 187.925 387.870 188.395 ;
        RECT 0.000 187.660 387.870 187.925 ;
        RECT 0.000 187.190 1.230 187.660 ;
        RECT 386.640 187.190 387.870 187.660 ;
        RECT 0.000 173.945 387.870 187.190 ;
        RECT 0.000 173.475 3.010 173.945 ;
        RECT 384.860 173.475 387.870 173.945 ;
        RECT 0.000 173.210 387.870 173.475 ;
        RECT 0.000 172.740 1.230 173.210 ;
        RECT 386.640 172.740 387.870 173.210 ;
        RECT 0.000 159.495 387.870 172.740 ;
        RECT 0.000 159.025 3.010 159.495 ;
        RECT 384.860 159.025 387.870 159.495 ;
        RECT 0.000 158.760 387.870 159.025 ;
        RECT 0.000 158.290 1.230 158.760 ;
        RECT 386.640 158.290 387.870 158.760 ;
        RECT 0.000 145.045 387.870 158.290 ;
        RECT 0.000 144.575 3.010 145.045 ;
        RECT 384.860 144.575 387.870 145.045 ;
        RECT 0.000 144.310 387.870 144.575 ;
        RECT 0.000 143.840 1.230 144.310 ;
        RECT 386.640 143.840 387.870 144.310 ;
        RECT 0.000 130.595 387.870 143.840 ;
        RECT 0.000 130.125 3.010 130.595 ;
        RECT 384.860 130.125 387.870 130.595 ;
        RECT 0.000 129.860 387.870 130.125 ;
        RECT 0.000 129.390 1.230 129.860 ;
        RECT 386.640 129.390 387.870 129.860 ;
        RECT 0.000 116.145 387.870 129.390 ;
        RECT 0.000 115.675 3.010 116.145 ;
        RECT 384.860 115.675 387.870 116.145 ;
        RECT 0.000 115.410 387.870 115.675 ;
        RECT 0.000 114.940 1.230 115.410 ;
        RECT 386.640 114.940 387.870 115.410 ;
        RECT 0.000 101.695 387.870 114.940 ;
        RECT 0.000 101.225 3.010 101.695 ;
        RECT 384.860 101.225 387.870 101.695 ;
        RECT 0.000 100.960 387.870 101.225 ;
        RECT 0.000 100.490 1.230 100.960 ;
        RECT 386.640 100.490 387.870 100.960 ;
        RECT 0.000 87.245 387.870 100.490 ;
        RECT 0.000 86.775 3.010 87.245 ;
        RECT 384.860 86.775 387.870 87.245 ;
        RECT 0.000 86.510 387.870 86.775 ;
        RECT 0.000 86.040 1.230 86.510 ;
        RECT 386.640 86.040 387.870 86.510 ;
        RECT 0.000 72.510 387.870 86.040 ;
        RECT 0.000 72.040 1.780 72.510 ;
        RECT 179.080 72.040 208.790 72.510 ;
        RECT 386.090 72.040 387.870 72.510 ;
        RECT 0.000 71.470 387.870 72.040 ;
        RECT 0.000 71.000 1.140 71.470 ;
        RECT 179.080 71.000 208.790 71.470 ;
        RECT 386.730 71.000 387.870 71.470 ;
        RECT 0.000 68.265 387.870 71.000 ;
        RECT 0.000 67.265 0.980 68.265 ;
        RECT 179.080 67.265 208.790 68.265 ;
        RECT 386.890 67.265 387.870 68.265 ;
        RECT 0.000 66.205 387.870 67.265 ;
        RECT 0.980 57.860 386.890 66.205 ;
        RECT 0.000 55.365 387.870 57.860 ;
        RECT 0.000 54.815 4.030 55.365 ;
        RECT 383.840 54.815 387.870 55.365 ;
        RECT 0.000 54.440 387.870 54.815 ;
        RECT 0.960 52.260 386.910 54.440 ;
        RECT 0.000 51.815 387.870 52.260 ;
        RECT 0.000 51.175 4.030 51.815 ;
        RECT 178.430 51.175 209.440 51.815 ;
        RECT 383.840 51.175 387.870 51.815 ;
        RECT 0.000 51.025 387.870 51.175 ;
        RECT 0.000 50.385 3.900 51.025 ;
        RECT 383.970 50.385 387.870 51.025 ;
        RECT 0.000 49.245 387.870 50.385 ;
        RECT 0.000 48.840 4.030 49.245 ;
        RECT 0.960 48.605 4.030 48.840 ;
        RECT 383.840 48.840 387.870 49.245 ;
        RECT 383.840 48.605 386.910 48.840 ;
        RECT 0.960 48.405 386.910 48.605 ;
        RECT 0.960 47.765 4.030 48.405 ;
        RECT 383.840 47.765 386.910 48.405 ;
        RECT 0.960 47.565 386.910 47.765 ;
        RECT 0.960 46.925 4.030 47.565 ;
        RECT 178.430 46.925 209.440 47.565 ;
        RECT 383.840 46.925 386.910 47.565 ;
        RECT 0.960 45.065 386.910 46.925 ;
        RECT 0.000 43.845 387.870 45.065 ;
        RECT 0.000 43.205 4.030 43.845 ;
        RECT 383.840 43.205 387.870 43.845 ;
        RECT 0.000 42.655 387.870 43.205 ;
        RECT 0.000 42.015 4.030 42.655 ;
        RECT 383.840 42.015 387.870 42.655 ;
        RECT 0.000 41.865 387.870 42.015 ;
        RECT 0.000 41.645 4.030 41.865 ;
        RECT 0.960 41.285 4.030 41.645 ;
        RECT 383.840 41.645 387.870 41.865 ;
        RECT 383.840 41.285 386.910 41.645 ;
        RECT 0.960 39.690 386.910 41.285 ;
        RECT 0.960 39.535 4.030 39.690 ;
        RECT 0.000 39.050 4.030 39.535 ;
        RECT 383.840 39.535 386.910 39.690 ;
        RECT 383.840 39.050 387.870 39.535 ;
        RECT 0.000 38.315 387.870 39.050 ;
        RECT 0.000 37.675 4.030 38.315 ;
        RECT 383.840 37.675 387.870 38.315 ;
        RECT 0.000 36.115 387.870 37.675 ;
        RECT 0.960 35.425 386.910 36.115 ;
        RECT 0.960 34.785 4.030 35.425 ;
        RECT 383.840 34.785 386.910 35.425 ;
        RECT 0.960 34.310 386.910 34.785 ;
        RECT 0.000 33.960 387.870 34.310 ;
        RECT 0.000 33.320 4.030 33.960 ;
        RECT 383.840 33.320 387.870 33.960 ;
        RECT 0.000 33.170 387.870 33.320 ;
        RECT 0.000 32.590 4.030 33.170 ;
        RECT 383.840 32.590 387.870 33.170 ;
        RECT 0.000 31.650 387.870 32.590 ;
        RECT 0.000 31.070 4.030 31.650 ;
        RECT 383.840 31.070 387.870 31.650 ;
        RECT 0.000 30.890 387.870 31.070 ;
        RECT 0.960 29.310 386.910 30.890 ;
        RECT 0.000 27.440 387.870 29.310 ;
        RECT 0.000 26.860 4.030 27.440 ;
        RECT 383.840 26.860 387.870 27.440 ;
        RECT 0.000 26.710 387.870 26.860 ;
        RECT 0.000 25.890 4.030 26.710 ;
        RECT 0.960 25.810 4.030 25.890 ;
        RECT 383.840 25.890 387.870 26.710 ;
        RECT 383.840 25.810 386.910 25.890 ;
        RECT 0.960 24.690 386.910 25.810 ;
        RECT 0.960 24.370 178.430 24.690 ;
        RECT 209.440 24.370 386.910 24.690 ;
        RECT 0.960 24.310 4.030 24.370 ;
        RECT 0.000 23.790 4.030 24.310 ;
        RECT 383.840 24.310 386.910 24.370 ;
        RECT 178.430 23.790 209.440 24.110 ;
        RECT 383.840 23.790 387.870 24.310 ;
        RECT 0.000 21.325 387.870 23.790 ;
        RECT 0.000 20.745 4.030 21.325 ;
        RECT 383.840 20.745 387.870 21.325 ;
        RECT 0.000 20.595 387.870 20.745 ;
        RECT 0.000 20.495 4.030 20.595 ;
        RECT 0.960 20.235 4.030 20.495 ;
        RECT 0.000 19.895 4.030 20.235 ;
        RECT 383.840 20.495 387.870 20.595 ;
        RECT 383.840 20.235 386.910 20.495 ;
        RECT 383.840 19.895 387.870 20.235 ;
        RECT 0.000 19.745 387.870 19.895 ;
        RECT 0.000 19.165 4.030 19.745 ;
        RECT 383.840 19.165 387.870 19.745 ;
        RECT 0.000 18.615 387.870 19.165 ;
        RECT 0.960 18.355 386.910 18.615 ;
        RECT 0.000 18.205 387.870 18.355 ;
        RECT 0.000 17.625 4.030 18.205 ;
        RECT 383.840 17.625 387.870 18.205 ;
        RECT 0.000 17.475 387.870 17.625 ;
        RECT 0.000 16.895 4.030 17.475 ;
        RECT 383.840 16.895 387.870 17.475 ;
        RECT 0.000 16.745 387.870 16.895 ;
        RECT 0.000 15.745 4.030 16.745 ;
        RECT 178.430 15.745 209.440 15.865 ;
        RECT 383.840 15.745 387.870 16.745 ;
        RECT 0.000 14.935 387.870 15.745 ;
        RECT 0.960 14.295 4.030 14.935 ;
        RECT 178.430 14.295 209.440 14.355 ;
        RECT 383.840 14.295 386.910 14.935 ;
        RECT 0.960 14.145 386.910 14.295 ;
        RECT 0.960 13.565 4.030 14.145 ;
        RECT 383.840 13.565 386.910 14.145 ;
        RECT 0.960 13.355 386.910 13.565 ;
        RECT 0.000 9.935 387.870 13.355 ;
        RECT 0.960 8.355 386.910 9.935 ;
        RECT 0.000 4.935 387.870 8.355 ;
        RECT 0.960 4.880 386.910 4.935 ;
        RECT 0.960 4.010 4.030 4.880 ;
        RECT 383.840 4.010 386.910 4.880 ;
        RECT 0.960 3.870 386.910 4.010 ;
        RECT 0.960 3.360 4.030 3.870 ;
        RECT 0.000 3.000 4.030 3.360 ;
        RECT 383.840 3.360 386.910 3.870 ;
        RECT 383.840 3.000 387.870 3.360 ;
  END
END CF_SRAM_1024x32
END LIBRARY

