magic
tech sky130A
magscale 1 2
timestamp 1758543462
<< viali >>
rect 65717 52649 65751 52683
rect 65993 52445 66027 52479
rect 65717 50269 65751 50303
rect 65717 49725 65751 49759
rect 65717 49181 65751 49215
rect 65717 47005 65751 47039
rect 65993 47005 66027 47039
rect 65717 43741 65751 43775
rect 68109 42721 68143 42755
rect 65717 42653 65751 42687
rect 68753 42653 68787 42687
rect 66729 41769 66763 41803
rect 67373 41565 67407 41599
rect 66453 40681 66487 40715
rect 67097 40477 67131 40511
rect 65717 39593 65751 39627
rect 66361 39389 66395 39423
rect 65717 38505 65751 38539
rect 66361 38301 66395 38335
rect 65717 37961 65751 37995
rect 66361 37757 66395 37791
rect 65717 36329 65751 36363
rect 66361 36125 66395 36159
rect 67005 35785 67039 35819
rect 65717 35649 65751 35683
rect 66637 35105 66671 35139
rect 65717 35037 65751 35071
rect 65717 34697 65751 34731
rect 66361 34493 66395 34527
rect 65717 34153 65751 34187
rect 66361 33949 66395 33983
rect 65717 33065 65751 33099
rect 66361 32861 66395 32895
rect 65717 31977 65751 32011
rect 66361 31773 66395 31807
rect 65717 30889 65751 30923
rect 66361 30685 66395 30719
rect 65717 29801 65751 29835
rect 66361 29597 66395 29631
rect 65717 28441 65751 28475
rect 67005 28373 67039 28407
rect 65717 28169 65751 28203
rect 66269 27965 66303 27999
rect 65717 27557 65751 27591
rect 66361 27421 66395 27455
rect 66637 27013 66671 27047
rect 65717 26945 65751 26979
rect 65717 26537 65751 26571
rect 66361 26333 66395 26367
rect 65717 25449 65751 25483
rect 66269 25245 66303 25279
rect 66085 24769 66119 24803
rect 66637 24701 66671 24735
rect 65717 24565 65751 24599
rect 65993 24565 66027 24599
rect 65901 24361 65935 24395
rect 66637 24361 66671 24395
rect 66453 24157 66487 24191
rect 67281 24157 67315 24191
rect 65809 24021 65843 24055
rect 65717 23817 65751 23851
rect 66453 23817 66487 23851
rect 67189 23817 67223 23851
rect 66269 23613 66303 23647
rect 67097 23613 67131 23647
rect 67741 23613 67775 23647
rect 65901 23273 65935 23307
rect 66637 23273 66671 23307
rect 66545 23069 66579 23103
rect 67189 23069 67223 23103
rect 65717 22933 65751 22967
rect 65717 22729 65751 22763
rect 66269 22525 66303 22559
rect 65717 7497 65751 7531
rect 69213 7497 69247 7531
rect 66545 7361 66579 7395
rect 66545 6953 66579 6987
rect 69213 6953 69247 6987
rect 66545 6409 66579 6443
rect 69213 6409 69247 6443
rect 50721 5865 50755 5899
rect 51457 5865 51491 5899
rect 52193 5865 52227 5899
rect 53297 5865 53331 5899
rect 55873 5865 55907 5899
rect 59185 5865 59219 5899
rect 59369 5865 59403 5899
rect 59553 5865 59587 5899
rect 59737 5865 59771 5899
rect 60657 5865 60691 5899
rect 60841 5865 60875 5899
rect 61025 5865 61059 5899
rect 61209 5865 61243 5899
rect 63601 5865 63635 5899
rect 63785 5865 63819 5899
rect 63969 5865 64003 5899
rect 66545 5865 66579 5899
rect 69213 5865 69247 5899
rect 42717 5797 42751 5831
rect 44741 5797 44775 5831
rect 54769 5797 54803 5831
rect 49617 5729 49651 5763
rect 57345 5729 57379 5763
rect 42533 5661 42567 5695
rect 44097 5661 44131 5695
rect 48973 5661 49007 5695
rect 50077 5661 50111 5695
rect 50813 5661 50847 5695
rect 51549 5661 51583 5695
rect 52653 5661 52687 5695
rect 53389 5661 53423 5695
rect 54125 5661 54159 5695
rect 55229 5661 55263 5695
rect 55965 5661 55999 5695
rect 56609 5661 56643 5695
rect 56701 5661 56735 5695
rect 43913 5593 43947 5627
rect 54033 5593 54067 5627
rect 48789 5525 48823 5559
rect 62129 5525 62163 5559
rect 62313 5525 62347 5559
rect 62497 5525 62531 5559
rect 62681 5525 62715 5559
rect 31033 5321 31067 5355
rect 49065 5321 49099 5355
rect 66545 5321 66579 5355
rect 69213 5321 69247 5355
rect 30113 5253 30147 5287
rect 30757 5253 30791 5287
rect 31125 5253 31159 5287
rect 47317 5253 47351 5287
rect 48145 5253 48179 5287
rect 62129 5253 62163 5287
rect 30389 5185 30423 5219
rect 31493 5185 31527 5219
rect 32505 5185 32539 5219
rect 32321 5117 32355 5151
rect 44649 5117 44683 5151
rect 44833 5117 44867 5151
rect 45569 5117 45603 5151
rect 47593 5117 47627 5151
rect 48237 5117 48271 5151
rect 48421 5117 48455 5151
rect 50537 5117 50571 5151
rect 54309 5117 54343 5151
rect 29929 5049 29963 5083
rect 45477 5049 45511 5083
rect 34713 4981 34747 5015
rect 35173 4981 35207 5015
rect 51181 4981 51215 5015
rect 54953 4981 54987 5015
rect 59185 4981 59219 5015
rect 60565 4981 60599 5015
rect 63601 4981 63635 5015
rect 30205 4777 30239 4811
rect 31585 4777 31619 4811
rect 35725 4777 35759 4811
rect 62129 4777 62163 4811
rect 66545 4777 66579 4811
rect 69213 4777 69247 4811
rect 34621 4709 34655 4743
rect 61209 4709 61243 4743
rect 63601 4709 63635 4743
rect 29837 4641 29871 4675
rect 30021 4641 30055 4675
rect 32597 4641 32631 4675
rect 34780 4641 34814 4675
rect 35265 4641 35299 4675
rect 46765 4641 46799 4675
rect 28917 4573 28951 4607
rect 29101 4573 29135 4607
rect 29285 4573 29319 4607
rect 29561 4573 29595 4607
rect 30941 4573 30975 4607
rect 32781 4573 32815 4607
rect 34253 4573 34287 4607
rect 34897 4573 34931 4607
rect 45569 4573 45603 4607
rect 47501 4573 47535 4607
rect 60565 4573 60599 4607
rect 28641 4505 28675 4539
rect 30481 4505 30515 4539
rect 30757 4505 30791 4539
rect 31426 4505 31460 4539
rect 33885 4505 33919 4539
rect 35449 4505 35483 4539
rect 48697 4505 48731 4539
rect 61050 4505 61084 4539
rect 29929 4437 29963 4471
rect 30665 4437 30699 4471
rect 31217 4437 31251 4471
rect 31309 4437 31343 4471
rect 32137 4437 32171 4471
rect 34989 4437 35023 4471
rect 59185 4437 59219 4471
rect 60841 4437 60875 4471
rect 60933 4437 60967 4471
rect 29745 4233 29779 4267
rect 30757 4233 30791 4267
rect 31585 4233 31619 4267
rect 32505 4233 32539 4267
rect 33701 4233 33735 4267
rect 33793 4233 33827 4267
rect 34345 4233 34379 4267
rect 34621 4233 34655 4267
rect 35081 4233 35115 4267
rect 35357 4233 35391 4267
rect 46949 4233 46983 4267
rect 48513 4233 48547 4267
rect 50169 4233 50203 4267
rect 51733 4233 51767 4267
rect 53205 4233 53239 4267
rect 54861 4233 54895 4267
rect 56333 4233 56367 4267
rect 58081 4233 58115 4267
rect 59369 4233 59403 4267
rect 60657 4233 60691 4267
rect 62313 4233 62347 4267
rect 63785 4233 63819 4267
rect 65257 4233 65291 4267
rect 66729 4233 66763 4267
rect 68385 4233 68419 4267
rect 69489 4233 69523 4267
rect 29377 4165 29411 4199
rect 29653 4165 29687 4199
rect 30849 4165 30883 4199
rect 32622 4165 32656 4199
rect 32965 4165 32999 4199
rect 34713 4165 34747 4199
rect 35240 4165 35274 4199
rect 35449 4165 35483 4199
rect 47041 4165 47075 4199
rect 48605 4165 48639 4199
rect 50261 4165 50295 4199
rect 51825 4165 51859 4199
rect 53297 4165 53331 4199
rect 54953 4165 54987 4199
rect 56425 4165 56459 4199
rect 58173 4165 58207 4199
rect 59461 4165 59495 4199
rect 62405 4165 62439 4199
rect 63877 4165 63911 4199
rect 63994 4165 64028 4199
rect 65349 4165 65383 4199
rect 66938 4165 66972 4199
rect 68477 4165 68511 4199
rect 69698 4165 69732 4199
rect 30297 4097 30331 4131
rect 31217 4097 31251 4131
rect 32137 4097 32171 4131
rect 35725 4097 35759 4131
rect 36001 4097 36035 4131
rect 36645 4097 36679 4131
rect 40693 4097 40727 4131
rect 47158 4097 47192 4131
rect 48237 4097 48271 4131
rect 49801 4097 49835 4131
rect 50378 4097 50412 4131
rect 51457 4097 51491 4131
rect 52929 4097 52963 4131
rect 54585 4097 54619 4131
rect 56057 4097 56091 4131
rect 57805 4097 57839 4131
rect 59093 4097 59127 4131
rect 62037 4097 62071 4131
rect 63509 4097 63543 4131
rect 65466 4097 65500 4131
rect 66821 4097 66855 4131
rect 68594 4097 68628 4131
rect 69581 4097 69615 4131
rect 28089 4029 28123 4063
rect 29193 4029 29227 4063
rect 29837 4029 29871 4063
rect 30389 4029 30423 4063
rect 30665 4029 30699 4063
rect 31493 4029 31527 4063
rect 31702 4029 31736 4063
rect 32413 4029 32447 4063
rect 33584 4029 33618 4063
rect 34069 4029 34103 4063
rect 34253 4029 34287 4063
rect 34504 4029 34538 4063
rect 34989 4029 35023 4063
rect 36277 4029 36311 4063
rect 40233 4029 40267 4063
rect 40785 4029 40819 4063
rect 46673 4029 46707 4063
rect 48722 4029 48756 4063
rect 49893 4029 49927 4063
rect 51365 4029 51399 4063
rect 51942 4029 51976 4063
rect 53414 4029 53448 4063
rect 54493 4029 54527 4063
rect 55070 4029 55104 4063
rect 55965 4029 55999 4063
rect 56542 4029 56576 4063
rect 58290 4029 58324 4063
rect 59578 4029 59612 4063
rect 62522 4029 62556 4063
rect 64981 4029 65015 4063
rect 66453 4029 66487 4063
rect 68109 4029 68143 4063
rect 69213 4029 69247 4063
rect 30021 3961 30055 3995
rect 35817 3961 35851 3995
rect 46581 3961 46615 3995
rect 47317 3961 47351 3995
rect 48881 3961 48915 3995
rect 50537 3961 50571 3995
rect 52101 3961 52135 3995
rect 55229 3961 55263 3995
rect 59737 3961 59771 3995
rect 68753 3961 68787 3995
rect 27537 3893 27571 3927
rect 28641 3893 28675 3927
rect 31033 3893 31067 3927
rect 31861 3893 31895 3927
rect 32781 3893 32815 3927
rect 33425 3893 33459 3927
rect 48145 3893 48179 3927
rect 53573 3893 53607 3927
rect 56701 3893 56735 3927
rect 58449 3893 58483 3927
rect 62681 3893 62715 3927
rect 64153 3893 64187 3927
rect 65625 3893 65659 3927
rect 67097 3893 67131 3927
rect 69857 3893 69891 3927
rect 32781 3689 32815 3723
rect 34437 3689 34471 3723
rect 35725 3689 35759 3723
rect 37933 3689 37967 3723
rect 64981 3689 65015 3723
rect 66545 3689 66579 3723
rect 68109 3689 68143 3723
rect 69213 3689 69247 3723
rect 31677 3621 31711 3655
rect 32413 3621 32447 3655
rect 34713 3621 34747 3655
rect 35541 3621 35575 3655
rect 46765 3621 46799 3655
rect 62129 3621 62163 3655
rect 63601 3621 63635 3655
rect 65717 3621 65751 3655
rect 26893 3553 26927 3587
rect 28641 3553 28675 3587
rect 30481 3553 30515 3587
rect 31309 3553 31343 3587
rect 31401 3553 31435 3587
rect 31518 3553 31552 3587
rect 32045 3553 32079 3587
rect 32873 3553 32907 3587
rect 34872 3553 34906 3587
rect 35357 3553 35391 3587
rect 36185 3553 36219 3587
rect 41337 3553 41371 3587
rect 64337 3553 64371 3587
rect 27077 3485 27111 3519
rect 27169 3485 27203 3519
rect 27997 3485 28031 3519
rect 29193 3485 29227 3519
rect 29469 3485 29503 3519
rect 30205 3485 30239 3519
rect 31033 3485 31067 3519
rect 31769 3485 31803 3519
rect 32254 3485 32288 3519
rect 32597 3485 32631 3519
rect 33149 3485 33183 3519
rect 33358 3485 33392 3519
rect 33609 3485 33643 3519
rect 35081 3485 35115 3519
rect 36369 3485 36403 3519
rect 36921 3485 36955 3519
rect 57621 3485 57655 3519
rect 63785 3485 63819 3519
rect 28549 3417 28583 3451
rect 29745 3417 29779 3451
rect 30113 3417 30147 3451
rect 30665 3417 30699 3451
rect 30941 3417 30975 3451
rect 34094 3417 34128 3451
rect 36553 3417 36587 3451
rect 38025 3417 38059 3451
rect 41613 3417 41647 3451
rect 58817 3417 58851 3451
rect 65901 3417 65935 3451
rect 27813 3349 27847 3383
rect 30573 3349 30607 3383
rect 32137 3349 32171 3383
rect 33241 3349 33275 3383
rect 33517 3349 33551 3383
rect 33885 3349 33919 3383
rect 33977 3349 34011 3383
rect 34253 3349 34287 3383
rect 34989 3349 35023 3383
rect 53021 3349 53055 3383
rect 59185 3349 59219 3383
rect 60565 3349 60599 3383
rect 28089 3145 28123 3179
rect 29561 3145 29595 3179
rect 31861 3145 31895 3179
rect 32781 3145 32815 3179
rect 33149 3145 33183 3179
rect 41981 3145 42015 3179
rect 44557 3145 44591 3179
rect 45385 3145 45419 3179
rect 57897 3145 57931 3179
rect 59093 3145 59127 3179
rect 59553 3145 59587 3179
rect 63509 3145 63543 3179
rect 66545 3145 66579 3179
rect 69213 3145 69247 3179
rect 26433 3077 26467 3111
rect 34713 3077 34747 3111
rect 60565 3077 60599 3111
rect 62129 3077 62163 3111
rect 25697 3009 25731 3043
rect 26709 3009 26743 3043
rect 27445 3009 27479 3043
rect 28733 3009 28767 3043
rect 31125 3009 31159 3043
rect 34989 3009 35023 3043
rect 37657 3009 37691 3043
rect 38393 3009 38427 3043
rect 38853 3009 38887 3043
rect 39129 3009 39163 3043
rect 41337 3009 41371 3043
rect 41613 3009 41647 3043
rect 42073 3009 42107 3043
rect 44649 3009 44683 3043
rect 45189 3009 45223 3043
rect 58173 3009 58207 3043
rect 59645 3009 59679 3043
rect 64613 3009 64647 3043
rect 69397 3009 69431 3043
rect 25973 2941 26007 2975
rect 28825 2941 28859 2975
rect 30113 2941 30147 2975
rect 30941 2941 30975 2975
rect 32229 2941 32263 2975
rect 36553 2941 36587 2975
rect 37473 2941 37507 2975
rect 37841 2941 37875 2975
rect 42349 2941 42383 2975
rect 44005 2941 44039 2975
rect 44925 2941 44959 2975
rect 63969 2941 64003 2975
rect 65073 2941 65107 2975
rect 67189 2941 67223 2975
rect 69857 2941 69891 2975
rect 29469 2873 29503 2907
rect 32965 2873 32999 2907
rect 35081 2873 35115 2907
rect 27997 2805 28031 2839
rect 30297 2805 30331 2839
rect 31217 2805 31251 2839
rect 33241 2805 33275 2839
rect 36001 2805 36035 2839
rect 42993 2805 43027 2839
rect 64521 2805 64555 2839
rect 67741 2805 67775 2839
rect 26709 2601 26743 2635
rect 29285 2601 29319 2635
rect 31401 2601 31435 2635
rect 33609 2601 33643 2635
rect 36645 2601 36679 2635
rect 37749 2601 37783 2635
rect 37841 2601 37875 2635
rect 39405 2601 39439 2635
rect 41613 2601 41647 2635
rect 41705 2601 41739 2635
rect 42441 2601 42475 2635
rect 44557 2601 44591 2635
rect 46029 2601 46063 2635
rect 52745 2601 52779 2635
rect 63509 2601 63543 2635
rect 66177 2601 66211 2635
rect 66545 2601 66579 2635
rect 69213 2601 69247 2635
rect 29653 2533 29687 2567
rect 48697 2533 48731 2567
rect 57345 2533 57379 2567
rect 25973 2465 26007 2499
rect 30573 2465 30607 2499
rect 34253 2465 34287 2499
rect 36001 2465 36035 2499
rect 42993 2465 43027 2499
rect 58081 2465 58115 2499
rect 59093 2465 59127 2499
rect 60565 2465 60599 2499
rect 64153 2465 64187 2499
rect 65533 2465 65567 2499
rect 67097 2465 67131 2499
rect 68385 2465 68419 2499
rect 71605 2465 71639 2499
rect 24961 2397 24995 2431
rect 26157 2397 26191 2431
rect 28181 2397 28215 2431
rect 28365 2397 28399 2431
rect 28733 2397 28767 2431
rect 30849 2397 30883 2431
rect 31493 2397 31527 2431
rect 32321 2397 32355 2431
rect 33057 2397 33091 2431
rect 33701 2397 33735 2431
rect 35633 2397 35667 2431
rect 37105 2397 37139 2431
rect 38393 2397 38427 2431
rect 38761 2397 38795 2431
rect 40601 2397 40635 2431
rect 41061 2397 41095 2431
rect 42349 2397 42383 2431
rect 43177 2397 43211 2431
rect 43821 2397 43855 2431
rect 43913 2397 43947 2431
rect 45201 2397 45235 2431
rect 45753 2397 45787 2431
rect 45845 2397 45879 2431
rect 46489 2397 46523 2431
rect 47501 2397 47535 2431
rect 48881 2397 48915 2431
rect 48973 2397 49007 2431
rect 49525 2397 49559 2431
rect 50169 2397 50203 2431
rect 51733 2397 51767 2431
rect 53665 2397 53699 2431
rect 55321 2397 55355 2431
rect 56333 2397 56367 2431
rect 57621 2397 57655 2431
rect 59277 2397 59311 2431
rect 61853 2397 61887 2431
rect 62313 2397 62347 2431
rect 63693 2397 63727 2431
rect 66637 2397 66671 2431
rect 68109 2397 68143 2431
rect 69489 2397 69523 2431
rect 70685 2397 70719 2431
rect 71329 2397 71363 2431
rect 71421 2397 71455 2431
rect 72617 2397 72651 2431
rect 26985 2329 27019 2363
rect 29837 2329 29871 2363
rect 30021 2329 30055 2363
rect 35081 2329 35115 2363
rect 40325 2329 40359 2363
rect 52285 2329 52319 2363
rect 52469 2329 52503 2363
rect 54217 2329 54251 2363
rect 54401 2329 54435 2363
rect 54769 2329 54803 2363
rect 56885 2329 56919 2363
rect 57069 2329 57103 2363
rect 61117 2329 61151 2363
rect 61301 2329 61335 2363
rect 72341 2329 72375 2363
rect 25145 2261 25179 2295
rect 25329 2261 25363 2295
rect 28457 2261 28491 2295
rect 32137 2261 32171 2295
rect 32873 2261 32907 2295
rect 47041 2261 47075 2295
rect 48145 2261 48179 2295
rect 50813 2261 50847 2295
rect 55873 2261 55907 2295
rect 59921 2261 59955 2295
rect 61025 2261 61059 2295
rect 62129 2261 62163 2295
rect 62865 2261 62899 2295
rect 70041 2261 70075 2295
rect 24409 2057 24443 2091
rect 25237 2057 25271 2091
rect 25973 2057 26007 2091
rect 26709 2057 26743 2091
rect 27077 2057 27111 2091
rect 36277 2057 36311 2091
rect 37013 2057 37047 2091
rect 40693 2057 40727 2091
rect 41429 2057 41463 2091
rect 45385 2057 45419 2091
rect 46949 2057 46983 2091
rect 47593 2057 47627 2091
rect 49433 2057 49467 2091
rect 50445 2057 50479 2091
rect 52653 2057 52687 2091
rect 55597 2057 55631 2091
rect 59093 2057 59127 2091
rect 59461 2057 59495 2091
rect 60565 2057 60599 2091
rect 61393 2057 61427 2091
rect 66545 2057 66579 2091
rect 69121 2057 69155 2091
rect 30205 1989 30239 2023
rect 62129 1989 62163 2023
rect 62589 1989 62623 2023
rect 67649 1989 67683 2023
rect 69213 1989 69247 2023
rect 71145 1989 71179 2023
rect 24225 1921 24259 1955
rect 26893 1921 26927 1955
rect 27445 1921 27479 1955
rect 29101 1921 29135 1955
rect 31861 1921 31895 1955
rect 33517 1921 33551 1955
rect 34161 1921 34195 1955
rect 37197 1921 37231 1955
rect 39037 1921 39071 1955
rect 39221 1921 39255 1955
rect 40509 1921 40543 1955
rect 41245 1921 41279 1955
rect 41981 1921 42015 1955
rect 42441 1921 42475 1955
rect 43913 1921 43947 1955
rect 47041 1921 47075 1955
rect 47777 1921 47811 1955
rect 47961 1921 47995 1955
rect 50537 1921 50571 1955
rect 50721 1921 50755 1955
rect 53481 1921 53515 1955
rect 55781 1921 55815 1955
rect 56241 1921 56275 1955
rect 57805 1921 57839 1955
rect 60013 1921 60047 1955
rect 63509 1921 63543 1955
rect 63693 1921 63727 1955
rect 67281 1921 67315 1955
rect 67373 1921 67407 1955
rect 69397 1921 69431 1955
rect 70869 1921 70903 1955
rect 71421 1921 71455 1955
rect 24593 1853 24627 1887
rect 25421 1853 25455 1887
rect 26157 1853 26191 1887
rect 28457 1853 28491 1887
rect 30665 1853 30699 1887
rect 32505 1853 32539 1887
rect 34713 1853 34747 1887
rect 35633 1853 35667 1887
rect 36461 1853 36495 1887
rect 37657 1853 37691 1887
rect 39865 1853 39899 1887
rect 39957 1853 39991 1887
rect 42901 1853 42935 1887
rect 44373 1853 44407 1887
rect 45937 1853 45971 1887
rect 46305 1853 46339 1887
rect 48421 1853 48455 1887
rect 49985 1853 50019 1887
rect 51181 1853 51215 1887
rect 53205 1853 53239 1887
rect 53941 1853 53975 1887
rect 54953 1853 54987 1887
rect 56701 1853 56735 1887
rect 60749 1853 60783 1887
rect 64153 1853 64187 1887
rect 65717 1853 65751 1887
rect 66361 1853 66395 1887
rect 66637 1853 66671 1887
rect 68569 1853 68603 1887
rect 69857 1853 69891 1887
rect 71881 1853 71915 1887
rect 38853 1785 38887 1819
rect 47225 1785 47259 1819
rect 56057 1785 56091 1819
rect 62405 1785 62439 1819
rect 58449 1717 58483 1751
rect 30389 1513 30423 1547
rect 35449 1513 35483 1547
rect 38117 1513 38151 1547
rect 41245 1513 41279 1547
rect 59093 1513 59127 1547
rect 66545 1513 66579 1547
rect 68293 1513 68327 1547
rect 69213 1513 69247 1547
rect 69581 1513 69615 1547
rect 60565 1445 60599 1479
rect 62129 1445 62163 1479
rect 63509 1445 63543 1479
rect 24501 1377 24535 1411
rect 46673 1377 46707 1411
rect 50537 1377 50571 1411
rect 71145 1377 71179 1411
rect 23581 1309 23615 1343
rect 25697 1309 25731 1343
rect 26157 1309 26191 1343
rect 26709 1309 26743 1343
rect 27261 1309 27295 1343
rect 29285 1309 29319 1343
rect 29837 1309 29871 1343
rect 30481 1309 30515 1343
rect 32045 1309 32079 1343
rect 32689 1309 32723 1343
rect 32781 1309 32815 1343
rect 33977 1309 34011 1343
rect 34897 1309 34931 1343
rect 35541 1309 35575 1343
rect 37565 1309 37599 1343
rect 38209 1309 38243 1343
rect 39773 1309 39807 1343
rect 41797 1309 41831 1343
rect 42349 1309 42383 1343
rect 43821 1309 43855 1343
rect 44373 1309 44407 1343
rect 45201 1309 45235 1343
rect 47225 1309 47259 1343
rect 47501 1309 47535 1343
rect 48973 1309 49007 1343
rect 49525 1309 49559 1343
rect 50077 1309 50111 1343
rect 52101 1309 52135 1343
rect 52653 1309 52687 1343
rect 54125 1309 54159 1343
rect 54677 1309 54711 1343
rect 55229 1309 55263 1343
rect 56701 1309 56735 1343
rect 57253 1309 57287 1343
rect 59277 1309 59311 1343
rect 59829 1309 59863 1343
rect 61301 1309 61335 1343
rect 61945 1309 61979 1343
rect 63693 1309 63727 1343
rect 66085 1309 66119 1343
rect 67005 1309 67039 1343
rect 67649 1309 67683 1343
rect 70133 1309 70167 1343
rect 70685 1309 70719 1343
rect 72157 1309 72191 1343
rect 72801 1309 72835 1343
rect 73813 1309 73847 1343
rect 28365 1241 28399 1275
rect 31677 1241 31711 1275
rect 36461 1241 36495 1275
rect 39129 1241 39163 1275
rect 40693 1241 40727 1275
rect 43269 1241 43303 1275
rect 46121 1241 46155 1275
rect 48421 1241 48455 1275
rect 53573 1241 53607 1275
rect 56149 1241 56183 1275
rect 64613 1241 64647 1275
rect 65533 1241 65567 1275
rect 68201 1241 68235 1275
rect 73261 1241 73295 1275
rect 23765 1173 23799 1207
rect 27813 1173 27847 1207
rect 51549 1173 51583 1207
<< metal1 >>
rect 65412 85978 74980 86000
rect 65412 85926 74210 85978
rect 74262 85926 74274 85978
rect 74326 85926 74338 85978
rect 74390 85926 74402 85978
rect 74454 85926 74466 85978
rect 74518 85926 74980 85978
rect 65412 85904 74980 85926
rect 65412 85434 74980 85456
rect 65412 85382 71858 85434
rect 71910 85382 71922 85434
rect 71974 85382 71986 85434
rect 72038 85382 72050 85434
rect 72102 85382 72114 85434
rect 72166 85382 74980 85434
rect 65412 85360 74980 85382
rect 65412 84890 74980 84912
rect 65412 84838 74210 84890
rect 74262 84838 74274 84890
rect 74326 84838 74338 84890
rect 74390 84838 74402 84890
rect 74454 84838 74466 84890
rect 74518 84838 74980 84890
rect 65412 84816 74980 84838
rect 65412 84346 74980 84368
rect 65412 84294 71858 84346
rect 71910 84294 71922 84346
rect 71974 84294 71986 84346
rect 72038 84294 72050 84346
rect 72102 84294 72114 84346
rect 72166 84294 74980 84346
rect 65412 84272 74980 84294
rect 63494 84232 63500 84244
rect 63328 84204 63500 84232
rect 63494 84192 63500 84204
rect 63552 84192 63558 84244
rect 65412 83802 74980 83824
rect 65412 83750 74210 83802
rect 74262 83750 74274 83802
rect 74326 83750 74338 83802
rect 74390 83750 74402 83802
rect 74454 83750 74466 83802
rect 74518 83750 74980 83802
rect 65412 83728 74980 83750
rect 65412 83258 74980 83280
rect 63328 83144 63356 83256
rect 65412 83206 71858 83258
rect 71910 83206 71922 83258
rect 71974 83206 71986 83258
rect 72038 83206 72050 83258
rect 72102 83206 72114 83258
rect 72166 83206 74980 83258
rect 65412 83184 74980 83206
rect 66898 83144 66904 83156
rect 63328 83116 66904 83144
rect 66898 83104 66904 83116
rect 66956 83104 66962 83156
rect 69198 83076 69204 83088
rect 63512 83048 69204 83076
rect 63512 83018 63540 83048
rect 69198 83036 69204 83048
rect 69256 83036 69262 83088
rect 63342 82990 63540 83018
rect 65412 82714 74980 82736
rect 65412 82662 74210 82714
rect 74262 82662 74274 82714
rect 74326 82662 74338 82714
rect 74390 82662 74402 82714
rect 74454 82662 74466 82714
rect 74518 82662 74980 82714
rect 65412 82640 74980 82662
rect 63494 82396 63500 82408
rect 63328 82368 63500 82396
rect 63328 82052 63356 82368
rect 63494 82356 63500 82368
rect 63552 82356 63558 82408
rect 65412 82170 74980 82192
rect 65412 82118 71858 82170
rect 71910 82118 71922 82170
rect 71974 82118 71986 82170
rect 72038 82118 72050 82170
rect 72102 82118 72114 82170
rect 72166 82118 74980 82170
rect 65412 82096 74980 82118
rect 65412 81626 74980 81648
rect 65412 81574 74210 81626
rect 74262 81574 74274 81626
rect 74326 81574 74338 81626
rect 74390 81574 74402 81626
rect 74454 81574 74466 81626
rect 74518 81574 74980 81626
rect 65412 81552 74980 81574
rect 65412 81082 74980 81104
rect 63328 80968 63356 81076
rect 65412 81030 71858 81082
rect 71910 81030 71922 81082
rect 71974 81030 71986 81082
rect 72038 81030 72050 81082
rect 72102 81030 72114 81082
rect 72166 81030 74980 81082
rect 65412 81008 74980 81030
rect 66714 80968 66720 80980
rect 63328 80940 66720 80968
rect 66714 80928 66720 80940
rect 66772 80928 66778 80980
rect 63328 80628 63356 80824
rect 66990 80628 66996 80640
rect 63328 80600 66996 80628
rect 66990 80588 66996 80600
rect 67048 80588 67054 80640
rect 65412 80538 74980 80560
rect 65412 80486 74210 80538
rect 74262 80486 74274 80538
rect 74326 80486 74338 80538
rect 74390 80486 74402 80538
rect 74454 80486 74466 80538
rect 74518 80486 74980 80538
rect 65412 80464 74980 80486
rect 63494 80016 63500 80028
rect 63328 79988 63500 80016
rect 63328 79872 63356 79988
rect 63494 79976 63500 79988
rect 63552 79976 63558 80028
rect 65412 79994 74980 80016
rect 65412 79942 71858 79994
rect 71910 79942 71922 79994
rect 71974 79942 71986 79994
rect 72038 79942 72050 79994
rect 72102 79942 72114 79994
rect 72166 79942 74980 79994
rect 65412 79920 74980 79942
rect 65412 79450 74980 79472
rect 65412 79398 74210 79450
rect 74262 79398 74274 79450
rect 74326 79398 74338 79450
rect 74390 79398 74402 79450
rect 74454 79398 74466 79450
rect 74518 79398 74980 79450
rect 65412 79376 74980 79398
rect 65412 78906 74980 78928
rect 63328 78724 63356 78896
rect 65412 78854 71858 78906
rect 71910 78854 71922 78906
rect 71974 78854 71986 78906
rect 72038 78854 72050 78906
rect 72102 78854 72114 78906
rect 72166 78854 74980 78906
rect 65412 78832 74980 78854
rect 65610 78724 65616 78736
rect 63328 78696 65616 78724
rect 65610 78684 65616 78696
rect 65668 78684 65674 78736
rect 63328 78452 63356 78644
rect 67082 78452 67088 78464
rect 63328 78424 67088 78452
rect 67082 78412 67088 78424
rect 67140 78412 67146 78464
rect 65412 78362 74980 78384
rect 65412 78310 74210 78362
rect 74262 78310 74274 78362
rect 74326 78310 74338 78362
rect 74390 78310 74402 78362
rect 74454 78310 74466 78362
rect 74518 78310 74980 78362
rect 65412 78288 74980 78310
rect 63494 78044 63500 78056
rect 63328 78016 63500 78044
rect 63328 77432 63356 78016
rect 63494 78004 63500 78016
rect 63552 78004 63558 78056
rect 65412 77818 74980 77840
rect 65412 77766 71858 77818
rect 71910 77766 71922 77818
rect 71974 77766 71986 77818
rect 72038 77766 72050 77818
rect 72102 77766 72114 77818
rect 72166 77766 74980 77818
rect 65412 77744 74980 77766
rect 63586 77432 63592 77444
rect 63328 77404 63592 77432
rect 63586 77392 63592 77404
rect 63644 77392 63650 77444
rect 65412 77274 74980 77296
rect 65412 77222 74210 77274
rect 74262 77222 74274 77274
rect 74326 77222 74338 77274
rect 74390 77222 74402 77274
rect 74454 77222 74466 77274
rect 74518 77222 74980 77274
rect 65412 77200 74980 77222
rect 63494 76730 63500 76742
rect 63342 76702 63500 76730
rect 63494 76690 63500 76702
rect 63552 76690 63558 76742
rect 65412 76730 74980 76752
rect 65412 76678 71858 76730
rect 71910 76678 71922 76730
rect 71974 76678 71986 76730
rect 72038 76678 72050 76730
rect 72102 76678 72114 76730
rect 72166 76678 74980 76730
rect 65412 76656 74980 76678
rect 63328 76140 63356 76464
rect 65412 76186 74980 76208
rect 63678 76140 63684 76152
rect 63328 76112 63684 76140
rect 63678 76100 63684 76112
rect 63736 76100 63742 76152
rect 65412 76134 74210 76186
rect 74262 76134 74274 76186
rect 74326 76134 74338 76186
rect 74390 76134 74402 76186
rect 74454 76134 74466 76186
rect 74518 76134 74980 76186
rect 65412 76112 74980 76134
rect 63586 75800 63592 75812
rect 63328 75772 63592 75800
rect 63328 75512 63356 75772
rect 63586 75760 63592 75772
rect 63644 75760 63650 75812
rect 65412 75642 74980 75664
rect 65412 75590 71858 75642
rect 71910 75590 71922 75642
rect 71974 75590 71986 75642
rect 72038 75590 72050 75642
rect 72102 75590 72114 75642
rect 72166 75590 74980 75642
rect 65412 75568 74980 75590
rect 65412 75098 74980 75120
rect 65412 75046 74210 75098
rect 74262 75046 74274 75098
rect 74326 75046 74338 75098
rect 74390 75046 74402 75098
rect 74454 75046 74466 75098
rect 74518 75046 74980 75098
rect 65412 75024 74980 75046
rect 63862 74576 63868 74588
rect 63328 74548 63868 74576
rect 63328 74536 63356 74548
rect 63862 74536 63868 74548
rect 63920 74536 63926 74588
rect 65412 74554 74980 74576
rect 65412 74502 71858 74554
rect 71910 74502 71922 74554
rect 71974 74502 71986 74554
rect 72038 74502 72050 74554
rect 72102 74502 72114 74554
rect 72166 74502 74980 74554
rect 65412 74480 74980 74502
rect 63328 73964 63356 74284
rect 65412 74010 74980 74032
rect 64138 73964 64144 73976
rect 63328 73936 64144 73964
rect 64138 73924 64144 73936
rect 64196 73924 64202 73976
rect 65412 73958 74210 74010
rect 74262 73958 74274 74010
rect 74326 73958 74338 74010
rect 74390 73958 74402 74010
rect 74454 73958 74466 74010
rect 74518 73958 74980 74010
rect 65412 73936 74980 73958
rect 65412 73466 74980 73488
rect 65412 73414 71858 73466
rect 71910 73414 71922 73466
rect 71974 73414 71986 73466
rect 72038 73414 72050 73466
rect 72102 73414 72114 73466
rect 72166 73414 74980 73466
rect 65412 73392 74980 73414
rect 63328 73216 63356 73332
rect 63586 73216 63592 73228
rect 63328 73188 63592 73216
rect 63586 73176 63592 73188
rect 63644 73176 63650 73228
rect 65412 72922 74980 72944
rect 65412 72870 74210 72922
rect 74262 72870 74274 72922
rect 74326 72870 74338 72922
rect 74390 72870 74402 72922
rect 74454 72870 74466 72922
rect 74518 72870 74980 72922
rect 65412 72848 74980 72870
rect 65412 72378 74980 72400
rect 63328 72196 63356 72356
rect 65412 72326 71858 72378
rect 71910 72326 71922 72378
rect 71974 72326 71986 72378
rect 72038 72326 72050 72378
rect 72102 72326 72114 72378
rect 72166 72326 74980 72378
rect 65412 72304 74980 72326
rect 65702 72196 65708 72208
rect 63328 72168 65708 72196
rect 65702 72156 65708 72168
rect 65760 72156 65766 72208
rect 69014 72128 69020 72140
rect 63328 72100 69020 72128
rect 69014 72088 69020 72100
rect 69072 72088 69078 72140
rect 65412 71834 74980 71856
rect 65412 71782 74210 71834
rect 74262 71782 74274 71834
rect 74326 71782 74338 71834
rect 74390 71782 74402 71834
rect 74454 71782 74466 71834
rect 74518 71782 74980 71834
rect 65412 71760 74980 71782
rect 63494 71612 63500 71664
rect 63552 71652 63558 71664
rect 66162 71652 66168 71664
rect 63552 71624 66168 71652
rect 63552 71612 63558 71624
rect 66162 71612 66168 71624
rect 66220 71612 66226 71664
rect 65610 71544 65616 71596
rect 65668 71584 65674 71596
rect 66346 71584 66352 71596
rect 65668 71556 66352 71584
rect 65668 71544 65674 71556
rect 66346 71544 66352 71556
rect 66404 71544 66410 71596
rect 63586 71448 63592 71460
rect 63328 71420 63592 71448
rect 63328 70836 63356 71420
rect 63586 71408 63592 71420
rect 63644 71408 63650 71460
rect 65412 71290 74980 71312
rect 65412 71238 71858 71290
rect 71910 71238 71922 71290
rect 71974 71238 71986 71290
rect 72038 71238 72050 71290
rect 72102 71238 72114 71290
rect 72166 71238 74980 71290
rect 65412 71216 74980 71238
rect 63494 70836 63500 70848
rect 63328 70808 63500 70836
rect 63494 70796 63500 70808
rect 63552 70796 63558 70848
rect 65412 70746 74980 70768
rect 65412 70694 74210 70746
rect 74262 70694 74274 70746
rect 74326 70694 74338 70746
rect 74390 70694 74402 70746
rect 74454 70694 74466 70746
rect 74518 70694 74980 70746
rect 65412 70672 74980 70694
rect 65412 70202 74980 70224
rect 63328 70020 63356 70176
rect 65412 70150 71858 70202
rect 71910 70150 71922 70202
rect 71974 70150 71986 70202
rect 72038 70150 72050 70202
rect 72102 70150 72114 70202
rect 72166 70150 74980 70202
rect 65412 70128 74980 70150
rect 65610 70020 65616 70032
rect 63328 69992 65616 70020
rect 65610 69980 65616 69992
rect 65668 69980 65674 70032
rect 63328 69612 63356 69924
rect 65412 69658 74980 69680
rect 63770 69612 63776 69624
rect 63328 69584 63776 69612
rect 63770 69572 63776 69584
rect 63828 69572 63834 69624
rect 65412 69606 74210 69658
rect 74262 69606 74274 69658
rect 74326 69606 74338 69658
rect 74390 69606 74402 69658
rect 74454 69606 74466 69658
rect 74518 69606 74980 69658
rect 65412 69584 74980 69606
rect 65412 69114 74980 69136
rect 65412 69062 71858 69114
rect 71910 69062 71922 69114
rect 71974 69062 71986 69114
rect 72038 69062 72050 69114
rect 72102 69062 72114 69114
rect 72166 69062 74980 69114
rect 65412 69040 74980 69062
rect 63494 69000 63500 69012
rect 63328 68972 63500 69000
rect 63328 68660 63356 68972
rect 63494 68960 63500 68972
rect 63552 68960 63558 69012
rect 66622 68660 66628 68672
rect 63328 68632 66628 68660
rect 66622 68620 66628 68632
rect 66680 68620 66686 68672
rect 65412 68570 74980 68592
rect 65412 68518 74210 68570
rect 74262 68518 74274 68570
rect 74326 68518 74338 68570
rect 74390 68518 74402 68570
rect 74454 68518 74466 68570
rect 74518 68518 74980 68570
rect 65412 68496 74980 68518
rect 65412 68026 74980 68048
rect 63328 67844 63356 67996
rect 65412 67974 71858 68026
rect 71910 67974 71922 68026
rect 71974 67974 71986 68026
rect 72038 67974 72050 68026
rect 72102 67974 72114 68026
rect 72166 67974 74980 68026
rect 65412 67952 74980 67974
rect 63328 67816 63448 67844
rect 63328 67640 63356 67744
rect 63420 67708 63448 67816
rect 63420 67680 64920 67708
rect 64782 67640 64788 67652
rect 63328 67612 64788 67640
rect 64782 67600 64788 67612
rect 64840 67600 64846 67652
rect 64892 67572 64920 67680
rect 65426 67572 65432 67584
rect 64892 67544 65432 67572
rect 65426 67532 65432 67544
rect 65484 67532 65490 67584
rect 65412 67482 74980 67504
rect 65412 67430 74210 67482
rect 74262 67430 74274 67482
rect 74326 67430 74338 67482
rect 74390 67430 74402 67482
rect 74454 67430 74466 67482
rect 74518 67430 74980 67482
rect 65412 67408 74980 67430
rect 65412 66938 74980 66960
rect 65412 66886 71858 66938
rect 71910 66886 71922 66938
rect 71974 66886 71986 66938
rect 72038 66886 72050 66938
rect 72102 66886 72114 66938
rect 72166 66886 74980 66938
rect 65412 66864 74980 66886
rect 63328 66484 63356 66792
rect 63586 66484 63592 66496
rect 63328 66456 63592 66484
rect 63586 66444 63592 66456
rect 63644 66444 63650 66496
rect 65412 66394 74980 66416
rect 65412 66342 74210 66394
rect 74262 66342 74274 66394
rect 74326 66342 74338 66394
rect 74390 66342 74402 66394
rect 74454 66342 74466 66394
rect 74518 66342 74980 66394
rect 65412 66320 74980 66342
rect 65412 65850 74980 65872
rect 63328 65668 63356 65816
rect 65412 65798 71858 65850
rect 71910 65798 71922 65850
rect 71974 65798 71986 65850
rect 72038 65798 72050 65850
rect 72102 65798 72114 65850
rect 72166 65798 74980 65850
rect 65412 65776 74980 65798
rect 65334 65668 65340 65680
rect 63328 65640 65340 65668
rect 65334 65628 65340 65640
rect 65392 65628 65398 65680
rect 63328 65260 63356 65564
rect 66990 65492 66996 65544
rect 67048 65532 67054 65544
rect 68094 65532 68100 65544
rect 67048 65504 68100 65532
rect 67048 65492 67054 65504
rect 68094 65492 68100 65504
rect 68152 65492 68158 65544
rect 65412 65306 74980 65328
rect 63494 65260 63500 65272
rect 63328 65232 63500 65260
rect 63494 65220 63500 65232
rect 63552 65220 63558 65272
rect 65412 65254 74210 65306
rect 74262 65254 74274 65306
rect 74326 65254 74338 65306
rect 74390 65254 74402 65306
rect 74454 65254 74466 65306
rect 74518 65254 74980 65306
rect 65412 65232 74980 65254
rect 63586 64852 63592 64864
rect 63328 64824 63592 64852
rect 63328 64308 63356 64824
rect 63586 64812 63592 64824
rect 63644 64812 63650 64864
rect 65412 64762 74980 64784
rect 63586 64676 63592 64728
rect 63644 64716 63650 64728
rect 63770 64716 63776 64728
rect 63644 64688 63776 64716
rect 63644 64676 63650 64688
rect 63770 64676 63776 64688
rect 63828 64676 63834 64728
rect 65412 64710 71858 64762
rect 71910 64710 71922 64762
rect 71974 64710 71986 64762
rect 72038 64710 72050 64762
rect 72102 64710 72114 64762
rect 72166 64710 74980 64762
rect 65412 64688 74980 64710
rect 63770 64308 63776 64320
rect 63328 64280 63776 64308
rect 63770 64268 63776 64280
rect 63828 64268 63834 64320
rect 65412 64218 74980 64240
rect 65412 64166 74210 64218
rect 74262 64166 74274 64218
rect 74326 64166 74338 64218
rect 74390 64166 74402 64218
rect 74454 64166 74466 64218
rect 74518 64166 74980 64218
rect 65412 64144 74980 64166
rect 65412 63674 74980 63696
rect 63328 63628 63356 63636
rect 63954 63628 63960 63640
rect 63328 63600 63960 63628
rect 63954 63588 63960 63600
rect 64012 63588 64018 63640
rect 65412 63622 71858 63674
rect 71910 63622 71922 63674
rect 71974 63622 71986 63674
rect 72038 63622 72050 63674
rect 72102 63622 72114 63674
rect 72166 63622 74980 63674
rect 65412 63600 74980 63622
rect 63328 63220 63356 63384
rect 63494 63220 63500 63232
rect 63328 63192 63500 63220
rect 63494 63180 63500 63192
rect 63552 63180 63558 63232
rect 65412 63130 74980 63152
rect 65412 63078 74210 63130
rect 74262 63078 74274 63130
rect 74326 63078 74338 63130
rect 74390 63078 74402 63130
rect 74454 63078 74466 63130
rect 74518 63078 74980 63130
rect 65412 63056 74980 63078
rect 65412 62586 74980 62608
rect 65412 62534 71858 62586
rect 71910 62534 71922 62586
rect 71974 62534 71986 62586
rect 72038 62534 72050 62586
rect 72102 62534 72114 62586
rect 72166 62534 74980 62586
rect 65412 62512 74980 62534
rect 63328 62132 63356 62432
rect 63770 62132 63776 62144
rect 63328 62104 63776 62132
rect 63770 62092 63776 62104
rect 63828 62092 63834 62144
rect 63954 62024 63960 62076
rect 64012 62064 64018 62076
rect 65242 62064 65248 62076
rect 64012 62036 65248 62064
rect 64012 62024 64018 62036
rect 65242 62024 65248 62036
rect 65300 62024 65306 62076
rect 65412 62042 74980 62064
rect 65412 61990 74210 62042
rect 74262 61990 74274 62042
rect 74326 61990 74338 62042
rect 74390 61990 74402 62042
rect 74454 61990 74466 62042
rect 74518 61990 74980 62042
rect 65412 61968 74980 61990
rect 65412 61498 74980 61520
rect 63328 61316 63356 61456
rect 65412 61446 71858 61498
rect 71910 61446 71922 61498
rect 71974 61446 71986 61498
rect 72038 61446 72050 61498
rect 72102 61446 72114 61498
rect 72166 61446 74980 61498
rect 65412 61424 74980 61446
rect 63954 61316 63960 61328
rect 63328 61288 63960 61316
rect 63954 61276 63960 61288
rect 64012 61276 64018 61328
rect 63328 61044 63356 61204
rect 63494 61044 63500 61056
rect 63328 61016 63500 61044
rect 63494 61004 63500 61016
rect 63552 61004 63558 61056
rect 65412 60954 74980 60976
rect 65412 60902 74210 60954
rect 74262 60902 74274 60954
rect 74326 60902 74338 60954
rect 74390 60902 74402 60954
rect 74454 60902 74466 60954
rect 74518 60902 74980 60954
rect 65412 60880 74980 60902
rect 65412 60410 74980 60432
rect 65412 60358 71858 60410
rect 71910 60358 71922 60410
rect 71974 60358 71986 60410
rect 72038 60358 72050 60410
rect 72102 60358 72114 60410
rect 72166 60358 74980 60410
rect 65412 60336 74980 60358
rect 63328 59956 63356 60252
rect 63770 59956 63776 59968
rect 63328 59928 63776 59956
rect 63770 59916 63776 59928
rect 63828 59916 63834 59968
rect 65412 59866 74980 59888
rect 65412 59814 74210 59866
rect 74262 59814 74274 59866
rect 74326 59814 74338 59866
rect 74390 59814 74402 59866
rect 74454 59814 74466 59866
rect 74518 59814 74980 59866
rect 65412 59792 74980 59814
rect 65412 59322 74980 59344
rect 63328 59140 63356 59276
rect 65412 59270 71858 59322
rect 71910 59270 71922 59322
rect 71974 59270 71986 59322
rect 72038 59270 72050 59322
rect 72102 59270 72114 59322
rect 72166 59270 74980 59322
rect 65412 59248 74980 59270
rect 65150 59140 65156 59152
rect 63328 59112 65156 59140
rect 65150 59100 65156 59112
rect 65208 59100 65214 59152
rect 63328 58732 63356 59024
rect 65412 58778 74980 58800
rect 63494 58732 63500 58744
rect 63328 58704 63500 58732
rect 63494 58692 63500 58704
rect 63552 58692 63558 58744
rect 65412 58726 74210 58778
rect 74262 58726 74274 58778
rect 74326 58726 74338 58778
rect 74390 58726 74402 58778
rect 74454 58726 74466 58778
rect 74518 58726 74980 58778
rect 65412 58704 74980 58726
rect 65412 58234 74980 58256
rect 65412 58182 71858 58234
rect 71910 58182 71922 58234
rect 71974 58182 71986 58234
rect 72038 58182 72050 58234
rect 72102 58182 72114 58234
rect 72166 58182 74980 58234
rect 65412 58160 74980 58182
rect 63328 57984 63356 58072
rect 63770 57984 63776 57996
rect 63328 57956 63776 57984
rect 63770 57944 63776 57956
rect 63828 57944 63834 57996
rect 65412 57690 74980 57712
rect 65412 57638 74210 57690
rect 74262 57638 74274 57690
rect 74326 57638 74338 57690
rect 74390 57638 74402 57690
rect 74454 57638 74466 57690
rect 74518 57638 74980 57690
rect 65412 57616 74980 57638
rect 65412 57146 74980 57168
rect 63328 56964 63356 57096
rect 65412 57094 71858 57146
rect 71910 57094 71922 57146
rect 71974 57094 71986 57146
rect 72038 57094 72050 57146
rect 72102 57094 72114 57146
rect 72166 57094 74980 57146
rect 65412 57072 74980 57094
rect 65058 56964 65064 56976
rect 63328 56936 65064 56964
rect 65058 56924 65064 56936
rect 65116 56924 65122 56976
rect 63328 56692 63356 56844
rect 63494 56692 63500 56704
rect 63328 56664 63500 56692
rect 63494 56652 63500 56664
rect 63552 56652 63558 56704
rect 65412 56602 74980 56624
rect 65412 56550 74210 56602
rect 74262 56550 74274 56602
rect 74326 56550 74338 56602
rect 74390 56550 74402 56602
rect 74454 56550 74466 56602
rect 74518 56550 74980 56602
rect 65412 56528 74980 56550
rect 65412 56058 74980 56080
rect 65412 56006 71858 56058
rect 71910 56006 71922 56058
rect 71974 56006 71986 56058
rect 72038 56006 72050 56058
rect 72102 56006 72114 56058
rect 72166 56006 74980 56058
rect 65412 55984 74980 56006
rect 63328 55604 63356 55892
rect 63770 55604 63776 55616
rect 63328 55576 63776 55604
rect 63770 55564 63776 55576
rect 63828 55564 63834 55616
rect 65412 55514 74980 55536
rect 65412 55462 74210 55514
rect 74262 55462 74274 55514
rect 74326 55462 74338 55514
rect 74390 55462 74402 55514
rect 74454 55462 74466 55514
rect 74518 55462 74980 55514
rect 65412 55440 74980 55462
rect 63954 55224 63960 55276
rect 64012 55264 64018 55276
rect 64966 55264 64972 55276
rect 64012 55236 64972 55264
rect 64012 55224 64018 55236
rect 64966 55224 64972 55236
rect 65024 55224 65030 55276
rect 65412 54970 74980 54992
rect 65412 54918 71858 54970
rect 71910 54918 71922 54970
rect 71974 54918 71986 54970
rect 72038 54918 72050 54970
rect 72102 54918 72114 54970
rect 72166 54918 74980 54970
rect 63328 54788 63356 54916
rect 65412 54896 74980 54918
rect 64046 54788 64052 54800
rect 63328 54760 64052 54788
rect 64046 54748 64052 54760
rect 64104 54748 64110 54800
rect 63236 54652 63264 54664
rect 63494 54652 63500 54664
rect 63236 54624 63500 54652
rect 63494 54612 63500 54624
rect 63552 54612 63558 54664
rect 65412 54426 74980 54448
rect 65412 54374 74210 54426
rect 74262 54374 74274 54426
rect 74326 54374 74338 54426
rect 74390 54374 74402 54426
rect 74454 54374 74466 54426
rect 74518 54374 74980 54426
rect 65412 54352 74980 54374
rect 65412 53882 74980 53904
rect 65412 53830 71858 53882
rect 71910 53830 71922 53882
rect 71974 53830 71986 53882
rect 72038 53830 72050 53882
rect 72102 53830 72114 53882
rect 72166 53830 74980 53882
rect 65412 53808 74980 53830
rect 63328 53564 63356 53712
rect 63770 53564 63776 53576
rect 63328 53536 63776 53564
rect 63770 53524 63776 53536
rect 63828 53524 63834 53576
rect 63328 53156 63356 53432
rect 65412 53338 74980 53360
rect 65412 53286 74210 53338
rect 74262 53286 74274 53338
rect 74326 53286 74338 53338
rect 74390 53286 74402 53338
rect 74454 53286 74466 53338
rect 74518 53286 74980 53338
rect 65412 53264 74980 53286
rect 66990 53156 66996 53168
rect 63328 53128 66996 53156
rect 66990 53116 66996 53128
rect 67048 53116 67054 53168
rect 65412 52794 74980 52816
rect 65412 52742 71858 52794
rect 71910 52742 71922 52794
rect 71974 52742 71986 52794
rect 72038 52742 72050 52794
rect 72102 52742 72114 52794
rect 72166 52742 74980 52794
rect 63328 52680 63356 52736
rect 65412 52720 74980 52742
rect 64690 52680 64696 52692
rect 63328 52652 64696 52680
rect 64690 52640 64696 52652
rect 64748 52640 64754 52692
rect 65705 52683 65763 52689
rect 65705 52680 65717 52683
rect 64846 52652 65717 52680
rect 63494 52572 63500 52624
rect 63552 52612 63558 52624
rect 64846 52612 64874 52652
rect 65705 52649 65717 52652
rect 65751 52649 65763 52683
rect 65705 52643 65763 52649
rect 69290 52612 69296 52624
rect 63552 52584 64874 52612
rect 64984 52584 69296 52612
rect 63552 52572 63558 52584
rect 64984 52544 65012 52584
rect 69290 52572 69296 52584
rect 69348 52572 69354 52624
rect 63696 52516 65012 52544
rect 63236 52476 63264 52484
rect 63696 52476 63724 52516
rect 65981 52479 66039 52485
rect 65981 52476 65993 52479
rect 63236 52448 63724 52476
rect 65260 52448 65993 52476
rect 65260 52408 65288 52448
rect 65981 52445 65993 52448
rect 66027 52445 66039 52479
rect 65981 52439 66039 52445
rect 63328 52380 65288 52408
rect 63328 52171 63356 52380
rect 65412 52250 74980 52272
rect 65412 52198 74210 52250
rect 74262 52198 74274 52250
rect 74326 52198 74338 52250
rect 74390 52198 74402 52250
rect 74454 52198 74466 52250
rect 74518 52198 74980 52250
rect 65412 52176 74980 52198
rect 63494 52108 63500 52120
rect 63342 52080 63500 52108
rect 63494 52068 63500 52080
rect 63552 52068 63558 52120
rect 65412 51706 74980 51728
rect 65412 51654 71858 51706
rect 71910 51654 71922 51706
rect 71974 51654 71986 51706
rect 72038 51654 72050 51706
rect 72102 51654 72114 51706
rect 72166 51654 74980 51706
rect 65412 51632 74980 51654
rect 63328 51524 63356 51532
rect 63770 51524 63776 51536
rect 63328 51496 63776 51524
rect 63770 51484 63776 51496
rect 63828 51524 63834 51536
rect 66530 51524 66536 51536
rect 63828 51496 66536 51524
rect 63828 51484 63834 51496
rect 66530 51484 66536 51496
rect 66588 51484 66594 51536
rect 65412 51162 74980 51184
rect 65412 51110 74210 51162
rect 74262 51110 74274 51162
rect 74326 51110 74338 51162
rect 74390 51110 74402 51162
rect 74454 51110 74466 51162
rect 74518 51110 74980 51162
rect 65412 51088 74980 51110
rect 65412 50618 74980 50640
rect 65412 50566 71858 50618
rect 71910 50566 71922 50618
rect 71974 50566 71986 50618
rect 72038 50566 72050 50618
rect 72102 50566 72114 50618
rect 72166 50566 74980 50618
rect 63328 50436 63356 50556
rect 65412 50544 74980 50566
rect 64874 50436 64880 50448
rect 63328 50408 64880 50436
rect 64874 50396 64880 50408
rect 64932 50396 64938 50448
rect 69106 50368 69112 50380
rect 64846 50340 69112 50368
rect 63236 50300 63264 50304
rect 64846 50300 64874 50340
rect 69106 50328 69112 50340
rect 69164 50328 69170 50380
rect 63236 50272 64874 50300
rect 65705 50303 65763 50309
rect 65705 50269 65717 50303
rect 65751 50269 65763 50303
rect 65705 50263 65763 50269
rect 65720 50232 65748 50263
rect 63328 50204 65748 50232
rect 63328 49996 63356 50204
rect 65412 50074 74980 50096
rect 65412 50022 74210 50074
rect 74262 50022 74274 50074
rect 74326 50022 74338 50074
rect 74390 50022 74402 50074
rect 74454 50022 74466 50074
rect 74518 50022 74980 50074
rect 65412 50000 74980 50022
rect 65705 49759 65763 49765
rect 65705 49756 65717 49759
rect 64846 49728 65717 49756
rect 64846 49688 64874 49728
rect 65705 49725 65717 49728
rect 65751 49725 65763 49759
rect 65705 49719 65763 49725
rect 63604 49671 64874 49688
rect 63342 49660 64874 49671
rect 63342 49643 63632 49660
rect 65412 49530 74980 49552
rect 65412 49478 71858 49530
rect 71910 49478 71922 49530
rect 71974 49478 71986 49530
rect 72038 49478 72050 49530
rect 72102 49478 72114 49530
rect 72166 49478 74980 49530
rect 65412 49456 74980 49478
rect 65705 49215 65763 49221
rect 65705 49212 65717 49215
rect 64846 49184 65717 49212
rect 63342 48804 63632 48809
rect 64322 48804 64328 48816
rect 63342 48781 64328 48804
rect 63604 48776 64328 48781
rect 64322 48764 64328 48776
rect 64380 48764 64386 48816
rect 64846 48736 64874 49184
rect 65705 49181 65717 49184
rect 65751 49181 65763 49215
rect 65705 49175 65763 49181
rect 65412 48986 74980 49008
rect 65412 48934 74210 48986
rect 74262 48934 74274 48986
rect 74326 48934 74338 48986
rect 74390 48934 74402 48986
rect 74454 48934 74466 48986
rect 74518 48934 74980 48986
rect 65412 48912 74980 48934
rect 63604 48729 64874 48736
rect 63342 48708 64874 48729
rect 63342 48701 63632 48708
rect 65412 48442 74980 48464
rect 65412 48390 71858 48442
rect 71910 48390 71922 48442
rect 71974 48390 71986 48442
rect 72038 48390 72050 48442
rect 72102 48390 72114 48442
rect 72166 48390 74980 48442
rect 65412 48368 74980 48390
rect 68554 48124 68560 48136
rect 63328 48096 68560 48124
rect 63328 48087 63356 48096
rect 68554 48084 68560 48096
rect 68612 48084 68618 48136
rect 63328 47716 63356 48007
rect 65412 47898 74980 47920
rect 65412 47846 74210 47898
rect 74262 47846 74274 47898
rect 74326 47846 74338 47898
rect 74390 47846 74402 47898
rect 74454 47846 74466 47898
rect 74518 47846 74980 47898
rect 65412 47824 74980 47846
rect 64414 47716 64420 47728
rect 63328 47688 64420 47716
rect 64414 47676 64420 47688
rect 64472 47676 64478 47728
rect 65518 47512 65524 47524
rect 63236 47484 65524 47512
rect 63236 47379 63264 47484
rect 65518 47472 65524 47484
rect 65576 47472 65582 47524
rect 65412 47354 74980 47376
rect 65412 47302 71858 47354
rect 71910 47302 71922 47354
rect 71974 47302 71986 47354
rect 72038 47302 72050 47354
rect 72102 47302 72114 47354
rect 72166 47302 74980 47354
rect 63328 47104 63356 47299
rect 65412 47280 74980 47302
rect 66070 47104 66076 47116
rect 63328 47076 66076 47104
rect 66070 47064 66076 47076
rect 66128 47064 66134 47116
rect 65702 46996 65708 47048
rect 65760 46996 65766 47048
rect 65978 46996 65984 47048
rect 66036 46996 66042 47048
rect 65412 46810 74980 46832
rect 65412 46758 74210 46810
rect 74262 46758 74274 46810
rect 74326 46758 74338 46810
rect 74390 46758 74402 46810
rect 74454 46758 74466 46810
rect 74518 46758 74980 46810
rect 65412 46736 74980 46758
rect 65412 46266 74980 46288
rect 65412 46214 71858 46266
rect 71910 46214 71922 46266
rect 71974 46214 71986 46266
rect 72038 46214 72050 46266
rect 72102 46214 72114 46266
rect 72166 46214 74980 46266
rect 65412 46192 74980 46214
rect 63342 45949 63632 45977
rect 63604 45948 63632 45949
rect 65794 45948 65800 45960
rect 63604 45920 65800 45948
rect 65794 45908 65800 45920
rect 65852 45908 65858 45960
rect 63328 45608 63356 45883
rect 65412 45722 74980 45744
rect 65412 45670 74210 45722
rect 74262 45670 74274 45722
rect 74326 45670 74338 45722
rect 74390 45670 74402 45722
rect 74454 45670 74466 45722
rect 74518 45670 74980 45722
rect 65412 45648 74980 45670
rect 65978 45608 65984 45620
rect 63328 45580 65984 45608
rect 65978 45568 65984 45580
rect 66036 45568 66042 45620
rect 63342 45268 63632 45269
rect 66438 45268 66444 45280
rect 63342 45241 66444 45268
rect 63604 45240 66444 45241
rect 66438 45228 66444 45240
rect 66496 45228 66502 45280
rect 65412 45178 74980 45200
rect 63328 44860 63356 45175
rect 65412 45126 71858 45178
rect 71910 45126 71922 45178
rect 71974 45126 71986 45178
rect 72038 45126 72050 45178
rect 72102 45126 72114 45178
rect 72166 45126 74980 45178
rect 65412 45104 74980 45126
rect 67174 44860 67180 44872
rect 63328 44832 67180 44860
rect 67174 44820 67180 44832
rect 67232 44820 67238 44872
rect 63678 44684 63684 44736
rect 63736 44724 63742 44736
rect 64230 44724 64236 44736
rect 63736 44696 64236 44724
rect 63736 44684 63742 44696
rect 64230 44684 64236 44696
rect 64288 44684 64294 44736
rect 65412 44634 74980 44656
rect 63678 44588 63684 44600
rect 63328 44560 63684 44588
rect 63328 44547 63356 44560
rect 63678 44548 63684 44560
rect 63736 44548 63742 44600
rect 65412 44582 74210 44634
rect 74262 44582 74274 44634
rect 74326 44582 74338 44634
rect 74390 44582 74402 44634
rect 74454 44582 74466 44634
rect 74518 44582 74980 44634
rect 65412 44560 74980 44582
rect 63328 44180 63356 44467
rect 67542 44180 67548 44192
rect 63328 44152 67548 44180
rect 67542 44140 67548 44152
rect 67600 44140 67606 44192
rect 65412 44090 74980 44112
rect 65412 44038 71858 44090
rect 71910 44038 71922 44090
rect 71974 44038 71986 44090
rect 72038 44038 72050 44090
rect 72102 44038 72114 44090
rect 72166 44038 74980 44090
rect 65412 44016 74980 44038
rect 64598 43840 64604 43852
rect 63328 43812 64604 43840
rect 64598 43800 64604 43812
rect 64656 43800 64662 43852
rect 65705 43775 65763 43781
rect 65705 43772 65717 43775
rect 63328 43744 65717 43772
rect 63328 43654 63356 43744
rect 65705 43741 65717 43744
rect 65751 43741 65763 43775
rect 65705 43735 65763 43741
rect 65518 43596 65524 43648
rect 65576 43636 65582 43648
rect 65886 43636 65892 43648
rect 65576 43608 65892 43636
rect 65576 43596 65582 43608
rect 65886 43596 65892 43608
rect 65944 43596 65950 43648
rect 65412 43546 74980 43568
rect 65412 43494 74210 43546
rect 74262 43494 74274 43546
rect 74326 43494 74338 43546
rect 74390 43494 74402 43546
rect 74454 43494 74466 43546
rect 74518 43494 74980 43546
rect 65412 43472 74980 43494
rect 64046 43392 64052 43444
rect 64104 43432 64110 43444
rect 65518 43432 65524 43444
rect 64104 43404 65524 43432
rect 64104 43392 64110 43404
rect 65518 43392 65524 43404
rect 65576 43392 65582 43444
rect 69382 43296 69388 43308
rect 63328 43268 69388 43296
rect 69382 43256 69388 43268
rect 69440 43256 69446 43308
rect 63328 42820 63356 43018
rect 65412 43002 74980 43024
rect 65412 42950 71858 43002
rect 71910 42950 71922 43002
rect 71974 42950 71986 43002
rect 72038 42950 72050 43002
rect 72102 42950 72114 43002
rect 72166 42950 74980 43002
rect 65412 42928 74980 42950
rect 63770 42820 63776 42832
rect 63328 42792 63776 42820
rect 63770 42780 63776 42792
rect 63828 42780 63834 42832
rect 66898 42712 66904 42764
rect 66956 42752 66962 42764
rect 68097 42755 68155 42761
rect 68097 42752 68109 42755
rect 66956 42724 68109 42752
rect 66956 42712 66962 42724
rect 68097 42721 68109 42724
rect 68143 42721 68155 42755
rect 68097 42715 68155 42721
rect 65705 42687 65763 42693
rect 65705 42684 65717 42687
rect 63328 42656 65717 42684
rect 63328 42402 63356 42656
rect 65705 42653 65717 42656
rect 65751 42653 65763 42687
rect 65705 42647 65763 42653
rect 68741 42687 68799 42693
rect 68741 42653 68753 42687
rect 68787 42684 68799 42687
rect 69658 42684 69664 42696
rect 68787 42656 69664 42684
rect 68787 42653 68799 42656
rect 68741 42647 68799 42653
rect 69658 42644 69664 42656
rect 69716 42644 69722 42696
rect 65412 42458 74980 42480
rect 65412 42406 74210 42458
rect 74262 42406 74274 42458
rect 74326 42406 74338 42458
rect 74390 42406 74402 42458
rect 74454 42406 74466 42458
rect 74518 42406 74980 42458
rect 65412 42384 74980 42406
rect 63328 41732 63356 42042
rect 65412 41914 74980 41936
rect 65412 41862 71858 41914
rect 71910 41862 71922 41914
rect 71974 41862 71986 41914
rect 72038 41862 72050 41914
rect 72102 41862 72114 41914
rect 72166 41862 74980 41914
rect 65412 41840 74980 41862
rect 66714 41760 66720 41812
rect 66772 41760 66778 41812
rect 63494 41732 63500 41744
rect 63328 41704 63500 41732
rect 63494 41692 63500 41704
rect 63552 41692 63558 41744
rect 67361 41599 67419 41605
rect 67361 41565 67373 41599
rect 67407 41596 67419 41599
rect 69842 41596 69848 41608
rect 67407 41568 69848 41596
rect 67407 41565 67419 41568
rect 67361 41559 67419 41565
rect 69842 41556 69848 41568
rect 69900 41556 69906 41608
rect 65412 41370 74980 41392
rect 65412 41318 74210 41370
rect 74262 41318 74274 41370
rect 74326 41318 74338 41370
rect 74390 41318 74402 41370
rect 74454 41318 74466 41370
rect 74518 41318 74980 41370
rect 65412 41296 74980 41318
rect 63328 40984 63356 41090
rect 63954 40984 63960 40996
rect 63328 40956 63960 40984
rect 63954 40944 63960 40956
rect 64012 40944 64018 40996
rect 65886 40876 65892 40928
rect 65944 40916 65950 40928
rect 66254 40916 66260 40928
rect 65944 40888 66260 40916
rect 65944 40876 65950 40888
rect 66254 40876 66260 40888
rect 66312 40876 66318 40928
rect 63328 40820 64874 40848
rect 64846 40644 64874 40820
rect 65412 40826 74980 40848
rect 65412 40774 71858 40826
rect 71910 40774 71922 40826
rect 71974 40774 71986 40826
rect 72038 40774 72050 40826
rect 72102 40774 72114 40826
rect 72166 40774 74980 40826
rect 65412 40752 74980 40774
rect 65886 40672 65892 40724
rect 65944 40712 65950 40724
rect 66070 40712 66076 40724
rect 65944 40684 66076 40712
rect 65944 40672 65950 40684
rect 66070 40672 66076 40684
rect 66128 40672 66134 40724
rect 66346 40672 66352 40724
rect 66404 40712 66410 40724
rect 66441 40715 66499 40721
rect 66441 40712 66453 40715
rect 66404 40684 66453 40712
rect 66404 40672 66410 40684
rect 66441 40681 66453 40684
rect 66487 40681 66499 40715
rect 66441 40675 66499 40681
rect 69474 40644 69480 40656
rect 64846 40616 69480 40644
rect 69474 40604 69480 40616
rect 69532 40604 69538 40656
rect 65518 40536 65524 40588
rect 65576 40576 65582 40588
rect 66070 40576 66076 40588
rect 65576 40548 66076 40576
rect 65576 40536 65582 40548
rect 66070 40536 66076 40548
rect 66128 40536 66134 40588
rect 67085 40511 67143 40517
rect 67085 40477 67097 40511
rect 67131 40508 67143 40511
rect 70026 40508 70032 40520
rect 67131 40480 70032 40508
rect 67131 40477 67143 40480
rect 67085 40471 67143 40477
rect 70026 40468 70032 40480
rect 70084 40468 70090 40520
rect 65412 40282 74980 40304
rect 65412 40230 74210 40282
rect 74262 40230 74274 40282
rect 74326 40230 74338 40282
rect 74390 40230 74402 40282
rect 74454 40230 74466 40282
rect 74518 40230 74980 40282
rect 65412 40208 74980 40230
rect 65058 40128 65064 40180
rect 65116 40168 65122 40180
rect 66346 40168 66352 40180
rect 65116 40140 66352 40168
rect 65116 40128 65122 40140
rect 66346 40128 66352 40140
rect 66404 40128 66410 40180
rect 64690 39992 64696 40044
rect 64748 40032 64754 40044
rect 65518 40032 65524 40044
rect 64748 40004 65524 40032
rect 64748 39992 64754 40004
rect 65518 39992 65524 40004
rect 65576 39992 65582 40044
rect 63328 39556 63356 39862
rect 65412 39738 74980 39760
rect 65412 39686 71858 39738
rect 71910 39686 71922 39738
rect 71974 39686 71986 39738
rect 72038 39686 72050 39738
rect 72102 39686 72114 39738
rect 72166 39686 74980 39738
rect 65412 39664 74980 39686
rect 65705 39627 65763 39633
rect 65705 39593 65717 39627
rect 65751 39624 65763 39627
rect 66162 39624 66168 39636
rect 65751 39596 66168 39624
rect 65751 39593 65763 39596
rect 65705 39587 65763 39593
rect 66162 39584 66168 39596
rect 66220 39584 66226 39636
rect 63494 39556 63500 39568
rect 63328 39528 63500 39556
rect 63494 39516 63500 39528
rect 63552 39516 63558 39568
rect 66349 39423 66407 39429
rect 66349 39389 66361 39423
rect 66395 39420 66407 39423
rect 68370 39420 68376 39432
rect 66395 39392 68376 39420
rect 66395 39389 66407 39392
rect 66349 39383 66407 39389
rect 68370 39380 68376 39392
rect 68428 39380 68434 39432
rect 65412 39194 74980 39216
rect 65412 39142 74210 39194
rect 74262 39142 74274 39194
rect 74326 39142 74338 39194
rect 74390 39142 74402 39194
rect 74454 39142 74466 39194
rect 74518 39142 74980 39194
rect 65412 39120 74980 39142
rect 63328 38740 63356 38910
rect 64046 38740 64052 38752
rect 63328 38712 64052 38740
rect 64046 38700 64052 38712
rect 64104 38700 64110 38752
rect 63862 38672 63868 38684
rect 63342 38644 63868 38672
rect 63862 38632 63868 38644
rect 63920 38632 63926 38684
rect 65412 38650 74980 38672
rect 65412 38598 71858 38650
rect 71910 38598 71922 38650
rect 71974 38598 71986 38650
rect 72038 38598 72050 38650
rect 72102 38598 72114 38650
rect 72166 38598 74980 38650
rect 65412 38576 74980 38598
rect 65702 38496 65708 38548
rect 65760 38496 65766 38548
rect 66349 38335 66407 38341
rect 66349 38301 66361 38335
rect 66395 38332 66407 38335
rect 68186 38332 68192 38344
rect 66395 38304 68192 38332
rect 66395 38301 66407 38304
rect 66349 38295 66407 38301
rect 68186 38292 68192 38304
rect 68244 38292 68250 38344
rect 65412 38106 74980 38128
rect 65412 38054 74210 38106
rect 74262 38054 74274 38106
rect 74326 38054 74338 38106
rect 74390 38054 74402 38106
rect 74454 38054 74466 38106
rect 74518 38054 74980 38106
rect 65412 38032 74980 38054
rect 63494 37992 63500 38004
rect 63328 37964 63500 37992
rect 63328 37380 63356 37964
rect 63494 37952 63500 37964
rect 63552 37952 63558 38004
rect 65610 37952 65616 38004
rect 65668 37992 65674 38004
rect 65705 37995 65763 38001
rect 65705 37992 65717 37995
rect 65668 37964 65717 37992
rect 65668 37952 65674 37964
rect 65705 37961 65717 37964
rect 65751 37961 65763 37995
rect 65705 37955 65763 37961
rect 63494 37816 63500 37868
rect 63552 37856 63558 37868
rect 63678 37856 63684 37868
rect 63552 37828 63684 37856
rect 63552 37816 63558 37828
rect 63678 37816 63684 37828
rect 63736 37816 63742 37868
rect 66349 37791 66407 37797
rect 66349 37757 66361 37791
rect 66395 37788 66407 37791
rect 66898 37788 66904 37800
rect 66395 37760 66904 37788
rect 66395 37757 66407 37760
rect 66349 37751 66407 37757
rect 66898 37748 66904 37760
rect 66956 37748 66962 37800
rect 65412 37562 74980 37584
rect 65412 37510 71858 37562
rect 71910 37510 71922 37562
rect 71974 37510 71986 37562
rect 72038 37510 72050 37562
rect 72102 37510 72114 37562
rect 72166 37510 74980 37562
rect 65412 37488 74980 37510
rect 63678 37380 63684 37392
rect 63328 37352 63684 37380
rect 63678 37340 63684 37352
rect 63736 37340 63742 37392
rect 65412 37018 74980 37040
rect 65412 36966 74210 37018
rect 74262 36966 74274 37018
rect 74326 36966 74338 37018
rect 74390 36966 74402 37018
rect 74454 36966 74466 37018
rect 74518 36966 74980 37018
rect 65412 36944 74980 36966
rect 63328 36564 63356 36730
rect 64506 36564 64512 36576
rect 63328 36536 64512 36564
rect 64506 36524 64512 36536
rect 64564 36524 64570 36576
rect 63328 36156 63356 36478
rect 65412 36474 74980 36496
rect 65412 36422 71858 36474
rect 71910 36422 71922 36474
rect 71974 36422 71986 36474
rect 72038 36422 72050 36474
rect 72102 36422 72114 36474
rect 72166 36422 74980 36474
rect 65412 36400 74980 36422
rect 65518 36320 65524 36372
rect 65576 36360 65582 36372
rect 65705 36363 65763 36369
rect 65705 36360 65717 36363
rect 65576 36332 65717 36360
rect 65576 36320 65582 36332
rect 65705 36329 65717 36332
rect 65751 36329 65763 36363
rect 65705 36323 65763 36329
rect 65426 36156 65432 36168
rect 63328 36128 65432 36156
rect 65426 36116 65432 36128
rect 65484 36116 65490 36168
rect 65518 36116 65524 36168
rect 65576 36156 65582 36168
rect 66070 36156 66076 36168
rect 65576 36128 66076 36156
rect 65576 36116 65582 36128
rect 66070 36116 66076 36128
rect 66128 36116 66134 36168
rect 66349 36159 66407 36165
rect 66349 36125 66361 36159
rect 66395 36156 66407 36159
rect 68278 36156 68284 36168
rect 66395 36128 68284 36156
rect 66395 36125 66407 36128
rect 66349 36119 66407 36125
rect 68278 36116 68284 36128
rect 68336 36116 68342 36168
rect 65412 35930 74980 35952
rect 65412 35878 74210 35930
rect 74262 35878 74274 35930
rect 74326 35878 74338 35930
rect 74390 35878 74402 35930
rect 74454 35878 74466 35930
rect 74518 35878 74980 35930
rect 65412 35856 74980 35878
rect 66990 35776 66996 35828
rect 67048 35776 67054 35828
rect 65702 35640 65708 35692
rect 65760 35640 65766 35692
rect 63328 35204 63356 35502
rect 65412 35386 74980 35408
rect 65412 35334 71858 35386
rect 71910 35334 71922 35386
rect 71974 35334 71986 35386
rect 72038 35334 72050 35386
rect 72102 35334 72114 35386
rect 72166 35334 74980 35386
rect 65412 35312 74980 35334
rect 63678 35204 63684 35216
rect 63328 35176 63684 35204
rect 63678 35164 63684 35176
rect 63736 35164 63742 35216
rect 65426 35204 65432 35216
rect 65260 35176 65432 35204
rect 65260 34660 65288 35176
rect 65426 35164 65432 35176
rect 65484 35164 65490 35216
rect 66622 35096 66628 35148
rect 66680 35096 66686 35148
rect 65426 35028 65432 35080
rect 65484 35068 65490 35080
rect 65705 35071 65763 35077
rect 65705 35068 65717 35071
rect 65484 35040 65717 35068
rect 65484 35028 65490 35040
rect 65705 35037 65717 35040
rect 65751 35037 65763 35071
rect 65705 35031 65763 35037
rect 65412 34842 74980 34864
rect 65412 34790 74210 34842
rect 74262 34790 74274 34842
rect 74326 34790 74338 34842
rect 74390 34790 74402 34842
rect 74454 34790 74466 34842
rect 74518 34790 74980 34842
rect 65412 34768 74980 34790
rect 65334 34688 65340 34740
rect 65392 34728 65398 34740
rect 65705 34731 65763 34737
rect 65705 34728 65717 34731
rect 65392 34700 65717 34728
rect 65392 34688 65398 34700
rect 65705 34697 65717 34700
rect 65751 34697 65763 34731
rect 65705 34691 65763 34697
rect 65260 34632 65380 34660
rect 65352 34604 65380 34632
rect 63328 34564 64874 34592
rect 63328 34550 63356 34564
rect 64846 34524 64874 34564
rect 65334 34552 65340 34604
rect 65392 34552 65398 34604
rect 67910 34592 67916 34604
rect 65444 34564 67916 34592
rect 65444 34524 65472 34564
rect 67910 34552 67916 34564
rect 67968 34552 67974 34604
rect 64846 34496 65472 34524
rect 66349 34527 66407 34533
rect 66349 34493 66361 34527
rect 66395 34524 66407 34527
rect 67358 34524 67364 34536
rect 66395 34496 67364 34524
rect 66395 34493 66407 34496
rect 66349 34487 66407 34493
rect 67358 34484 67364 34496
rect 67416 34484 67422 34536
rect 65412 34298 74980 34320
rect 63328 33980 63356 34298
rect 65412 34246 71858 34298
rect 71910 34246 71922 34298
rect 71974 34246 71986 34298
rect 72038 34246 72050 34298
rect 72102 34246 72114 34298
rect 72166 34246 74980 34298
rect 65412 34224 74980 34246
rect 65242 34144 65248 34196
rect 65300 34184 65306 34196
rect 65705 34187 65763 34193
rect 65705 34184 65717 34187
rect 65300 34156 65717 34184
rect 65300 34144 65306 34156
rect 65705 34153 65717 34156
rect 65751 34153 65763 34187
rect 65705 34147 65763 34153
rect 64690 33980 64696 33992
rect 63328 33952 64696 33980
rect 64690 33940 64696 33952
rect 64748 33940 64754 33992
rect 66349 33983 66407 33989
rect 66349 33949 66361 33983
rect 66395 33980 66407 33983
rect 67450 33980 67456 33992
rect 66395 33952 67456 33980
rect 66395 33949 66407 33952
rect 66349 33943 66407 33949
rect 67450 33940 67456 33952
rect 67508 33940 67514 33992
rect 65412 33754 74980 33776
rect 65412 33702 74210 33754
rect 74262 33702 74274 33754
rect 74326 33702 74338 33754
rect 74390 33702 74402 33754
rect 74454 33702 74466 33754
rect 74518 33702 74980 33754
rect 65412 33680 74980 33702
rect 63328 33164 63356 33322
rect 65412 33210 74980 33232
rect 63678 33164 63684 33176
rect 63328 33136 63684 33164
rect 63678 33124 63684 33136
rect 63736 33124 63742 33176
rect 65412 33158 71858 33210
rect 71910 33158 71922 33210
rect 71974 33158 71986 33210
rect 72038 33158 72050 33210
rect 72102 33158 72114 33210
rect 72166 33158 74980 33210
rect 65412 33136 74980 33158
rect 65150 33056 65156 33108
rect 65208 33096 65214 33108
rect 65705 33099 65763 33105
rect 65705 33096 65717 33099
rect 65208 33068 65717 33096
rect 65208 33056 65214 33068
rect 65705 33065 65717 33068
rect 65751 33065 65763 33099
rect 65705 33059 65763 33065
rect 66349 32895 66407 32901
rect 66349 32861 66361 32895
rect 66395 32892 66407 32895
rect 66622 32892 66628 32904
rect 66395 32864 66628 32892
rect 66395 32861 66407 32864
rect 66349 32855 66407 32861
rect 66622 32852 66628 32864
rect 66680 32852 66686 32904
rect 65412 32666 74980 32688
rect 65412 32614 74210 32666
rect 74262 32614 74274 32666
rect 74326 32614 74338 32666
rect 74390 32614 74402 32666
rect 74454 32614 74466 32666
rect 74518 32614 74980 32666
rect 65412 32592 74980 32614
rect 69566 32416 69572 32428
rect 63328 32388 69572 32416
rect 63328 32370 63356 32388
rect 69566 32376 69572 32388
rect 69624 32376 69630 32428
rect 65412 32122 74980 32144
rect 63328 31804 63356 32118
rect 65412 32070 71858 32122
rect 71910 32070 71922 32122
rect 71974 32070 71986 32122
rect 72038 32070 72050 32122
rect 72102 32070 72114 32122
rect 72166 32070 74980 32122
rect 65412 32048 74980 32070
rect 64966 31968 64972 32020
rect 65024 32008 65030 32020
rect 65705 32011 65763 32017
rect 65705 32008 65717 32011
rect 65024 31980 65717 32008
rect 65024 31968 65030 31980
rect 65705 31977 65717 31980
rect 65751 31977 65763 32011
rect 65705 31971 65763 31977
rect 66349 31807 66407 31813
rect 63328 31776 64184 31804
rect 64156 31668 64184 31776
rect 66349 31773 66361 31807
rect 66395 31804 66407 31807
rect 66806 31804 66812 31816
rect 66395 31776 66812 31804
rect 66395 31773 66407 31776
rect 66349 31767 66407 31773
rect 64230 31696 64236 31748
rect 64288 31736 64294 31748
rect 64288 31708 64460 31736
rect 64288 31696 64294 31708
rect 64156 31640 64276 31668
rect 63678 31600 63684 31612
rect 63328 31572 63684 31600
rect 63328 30852 63356 31572
rect 63678 31560 63684 31572
rect 63736 31560 63742 31612
rect 64248 31544 64276 31640
rect 64432 31544 64460 31708
rect 64506 31696 64512 31748
rect 64564 31696 64570 31748
rect 64598 31714 64604 31766
rect 64656 31714 64662 31766
rect 66806 31764 66812 31776
rect 66864 31764 66870 31816
rect 64524 31544 64552 31696
rect 64230 31492 64236 31544
rect 64288 31492 64294 31544
rect 64414 31492 64420 31544
rect 64472 31492 64478 31544
rect 64506 31492 64512 31544
rect 64564 31492 64570 31544
rect 63678 31424 63684 31476
rect 63736 31464 63742 31476
rect 64616 31464 64644 31714
rect 65412 31578 74980 31600
rect 65412 31526 74210 31578
rect 74262 31526 74274 31578
rect 74326 31526 74338 31578
rect 74390 31526 74402 31578
rect 74454 31526 74466 31578
rect 74518 31526 74980 31578
rect 65412 31504 74980 31526
rect 63736 31436 64644 31464
rect 63736 31424 63742 31436
rect 65412 31034 74980 31056
rect 65412 30982 71858 31034
rect 71910 30982 71922 31034
rect 71974 30982 71986 31034
rect 72038 30982 72050 31034
rect 72102 30982 72114 31034
rect 72166 30982 74980 31034
rect 65412 30960 74980 30982
rect 65058 30880 65064 30932
rect 65116 30920 65122 30932
rect 65705 30923 65763 30929
rect 65705 30920 65717 30923
rect 65116 30892 65717 30920
rect 65116 30880 65122 30892
rect 65705 30889 65717 30892
rect 65751 30889 65763 30923
rect 65705 30883 65763 30889
rect 65150 30852 65156 30864
rect 63328 30824 65156 30852
rect 65150 30812 65156 30824
rect 65208 30812 65214 30864
rect 66349 30719 66407 30725
rect 66349 30685 66361 30719
rect 66395 30716 66407 30719
rect 66714 30716 66720 30728
rect 66395 30688 66720 30716
rect 66395 30685 66407 30688
rect 66349 30679 66407 30685
rect 66714 30676 66720 30688
rect 66772 30676 66778 30728
rect 65412 30490 74980 30512
rect 65412 30438 74210 30490
rect 74262 30438 74274 30490
rect 74326 30438 74338 30490
rect 74390 30438 74402 30490
rect 74454 30438 74466 30490
rect 74518 30438 74980 30490
rect 65412 30416 74980 30438
rect 64414 30336 64420 30388
rect 64472 30376 64478 30388
rect 64966 30376 64972 30388
rect 64472 30348 64972 30376
rect 64472 30336 64478 30348
rect 64966 30336 64972 30348
rect 65024 30336 65030 30388
rect 63328 30172 63356 30190
rect 68002 30172 68008 30184
rect 63328 30144 68008 30172
rect 68002 30132 68008 30144
rect 68060 30132 68066 30184
rect 65412 29946 74980 29968
rect 63328 29764 63356 29938
rect 65412 29894 71858 29946
rect 71910 29894 71922 29946
rect 71974 29894 71986 29946
rect 72038 29894 72050 29946
rect 72102 29894 72114 29946
rect 72166 29894 74980 29946
rect 65412 29872 74980 29894
rect 65705 29835 65763 29841
rect 65705 29801 65717 29835
rect 65751 29832 65763 29835
rect 66162 29832 66168 29844
rect 65751 29804 66168 29832
rect 65751 29801 65763 29804
rect 65705 29795 65763 29801
rect 66162 29792 66168 29804
rect 66220 29792 66226 29844
rect 68462 29764 68468 29776
rect 63328 29736 68468 29764
rect 68462 29724 68468 29736
rect 68520 29724 68526 29776
rect 66346 29588 66352 29640
rect 66404 29588 66410 29640
rect 65412 29402 74980 29424
rect 65412 29350 74210 29402
rect 74262 29350 74274 29402
rect 74326 29350 74338 29402
rect 74390 29350 74402 29402
rect 74454 29350 74466 29402
rect 74518 29350 74980 29402
rect 65412 29328 74980 29350
rect 63328 28676 63356 28962
rect 65412 28858 74980 28880
rect 65412 28806 71858 28858
rect 71910 28806 71922 28858
rect 71974 28806 71986 28858
rect 72038 28806 72050 28858
rect 72102 28806 72114 28858
rect 72166 28806 74980 28858
rect 65412 28784 74980 28806
rect 65150 28676 65156 28688
rect 63328 28648 65156 28676
rect 65150 28636 65156 28648
rect 65208 28636 65214 28688
rect 65702 28432 65708 28484
rect 65760 28432 65766 28484
rect 65518 28364 65524 28416
rect 65576 28404 65582 28416
rect 66993 28407 67051 28413
rect 66993 28404 67005 28407
rect 65576 28376 67005 28404
rect 65576 28364 65582 28376
rect 66993 28373 67005 28376
rect 67039 28373 67051 28407
rect 66993 28367 67051 28373
rect 65412 28314 74980 28336
rect 65412 28262 74210 28314
rect 74262 28262 74274 28314
rect 74326 28262 74338 28314
rect 74390 28262 74402 28314
rect 74454 28262 74466 28314
rect 74518 28262 74980 28314
rect 65412 28240 74980 28262
rect 65334 28160 65340 28212
rect 65392 28200 65398 28212
rect 65705 28203 65763 28209
rect 65705 28200 65717 28203
rect 65392 28172 65717 28200
rect 65392 28160 65398 28172
rect 65705 28169 65717 28172
rect 65751 28169 65763 28203
rect 65705 28163 65763 28169
rect 63328 27928 63356 28010
rect 66254 27956 66260 28008
rect 66312 27956 66318 28008
rect 64414 27928 64420 27940
rect 63328 27900 64420 27928
rect 64414 27888 64420 27900
rect 64472 27888 64478 27940
rect 70118 27860 70124 27872
rect 63512 27832 70124 27860
rect 63512 27792 63540 27832
rect 70118 27820 70124 27832
rect 70176 27820 70182 27872
rect 63236 27764 63540 27792
rect 65412 27770 74980 27792
rect 63236 27758 63264 27764
rect 65412 27718 71858 27770
rect 71910 27718 71922 27770
rect 71974 27718 71986 27770
rect 72038 27718 72050 27770
rect 72102 27718 72114 27770
rect 72166 27718 74980 27770
rect 65412 27696 74980 27718
rect 65426 27548 65432 27600
rect 65484 27588 65490 27600
rect 65705 27591 65763 27597
rect 65705 27588 65717 27591
rect 65484 27560 65717 27588
rect 65484 27548 65490 27560
rect 65705 27557 65717 27560
rect 65751 27557 65763 27591
rect 65705 27551 65763 27557
rect 66349 27455 66407 27461
rect 66349 27421 66361 27455
rect 66395 27452 66407 27455
rect 67266 27452 67272 27464
rect 66395 27424 67272 27452
rect 66395 27421 66407 27424
rect 66349 27415 66407 27421
rect 67266 27412 67272 27424
rect 67324 27412 67330 27464
rect 65412 27226 74980 27248
rect 65412 27174 74210 27226
rect 74262 27174 74274 27226
rect 74326 27174 74338 27226
rect 74390 27174 74402 27226
rect 74454 27174 74466 27226
rect 74518 27174 74980 27226
rect 65412 27152 74980 27174
rect 66530 27004 66536 27056
rect 66588 27044 66594 27056
rect 66625 27047 66683 27053
rect 66625 27044 66637 27047
rect 66588 27016 66637 27044
rect 66588 27004 66594 27016
rect 66625 27013 66637 27016
rect 66671 27013 66683 27047
rect 66625 27007 66683 27013
rect 65610 26936 65616 26988
rect 65668 26976 65674 26988
rect 65705 26979 65763 26985
rect 65705 26976 65717 26979
rect 65668 26948 65717 26976
rect 65668 26936 65674 26948
rect 65705 26945 65717 26948
rect 65751 26945 65763 26979
rect 65705 26939 65763 26945
rect 63328 26772 63356 26782
rect 65150 26772 65156 26784
rect 63328 26744 65156 26772
rect 65150 26732 65156 26744
rect 65208 26732 65214 26784
rect 66622 26732 66628 26784
rect 66680 26772 66686 26784
rect 66806 26772 66812 26784
rect 66680 26744 66812 26772
rect 66680 26732 66686 26744
rect 66806 26732 66812 26744
rect 66864 26732 66870 26784
rect 65412 26682 74980 26704
rect 65412 26630 71858 26682
rect 71910 26630 71922 26682
rect 71974 26630 71986 26682
rect 72038 26630 72050 26682
rect 72102 26630 72114 26682
rect 72166 26630 74980 26682
rect 65412 26608 74980 26630
rect 64874 26528 64880 26580
rect 64932 26568 64938 26580
rect 65705 26571 65763 26577
rect 65705 26568 65717 26571
rect 64932 26540 65717 26568
rect 64932 26528 64938 26540
rect 65705 26537 65717 26540
rect 65751 26537 65763 26571
rect 65705 26531 65763 26537
rect 66349 26367 66407 26373
rect 66349 26333 66361 26367
rect 66395 26364 66407 26367
rect 66714 26364 66720 26376
rect 66395 26336 66720 26364
rect 66395 26333 66407 26336
rect 66349 26327 66407 26333
rect 66714 26324 66720 26336
rect 66772 26324 66778 26376
rect 65412 26138 74980 26160
rect 65412 26086 74210 26138
rect 74262 26086 74274 26138
rect 74326 26086 74338 26138
rect 74390 26086 74402 26138
rect 74454 26086 74466 26138
rect 74518 26086 74980 26138
rect 65412 26064 74980 26086
rect 63328 25684 63356 25830
rect 69934 25684 69940 25696
rect 63328 25656 69940 25684
rect 69934 25644 69940 25656
rect 69992 25644 69998 25696
rect 65412 25594 74980 25616
rect 63328 25276 63356 25578
rect 65412 25542 71858 25594
rect 71910 25542 71922 25594
rect 71974 25542 71986 25594
rect 72038 25542 72050 25594
rect 72102 25542 72114 25594
rect 72166 25542 74980 25594
rect 65412 25520 74980 25542
rect 64598 25440 64604 25492
rect 64656 25480 64662 25492
rect 65705 25483 65763 25489
rect 65705 25480 65717 25483
rect 64656 25452 65717 25480
rect 64656 25440 64662 25452
rect 65705 25449 65717 25452
rect 65751 25449 65763 25483
rect 65705 25443 65763 25449
rect 64598 25276 64604 25288
rect 63328 25248 64604 25276
rect 64598 25236 64604 25248
rect 64656 25236 64662 25288
rect 65426 25236 65432 25288
rect 65484 25276 65490 25288
rect 66257 25279 66315 25285
rect 66257 25276 66269 25279
rect 65484 25248 66269 25276
rect 65484 25236 65490 25248
rect 66257 25245 66269 25248
rect 66303 25245 66315 25279
rect 66257 25239 66315 25245
rect 65412 25050 74980 25072
rect 65412 24998 74210 25050
rect 74262 24998 74274 25050
rect 74326 24998 74338 25050
rect 74390 24998 74402 25050
rect 74454 24998 74466 25050
rect 74518 24998 74980 25050
rect 65412 24976 74980 24998
rect 66070 24760 66076 24812
rect 66128 24760 66134 24812
rect 66162 24692 66168 24744
rect 66220 24732 66226 24744
rect 66625 24735 66683 24741
rect 66625 24732 66637 24735
rect 66220 24704 66637 24732
rect 66220 24692 66226 24704
rect 66625 24701 66637 24704
rect 66671 24701 66683 24735
rect 66625 24695 66683 24701
rect 63328 24324 63356 24602
rect 65426 24556 65432 24608
rect 65484 24596 65490 24608
rect 65705 24599 65763 24605
rect 65705 24596 65717 24599
rect 65484 24568 65717 24596
rect 65484 24556 65490 24568
rect 65705 24565 65717 24568
rect 65751 24565 65763 24599
rect 65705 24559 65763 24565
rect 65981 24599 66039 24605
rect 65981 24565 65993 24599
rect 66027 24596 66039 24599
rect 66070 24596 66076 24608
rect 66027 24568 66076 24596
rect 66027 24565 66039 24568
rect 65981 24559 66039 24565
rect 66070 24556 66076 24568
rect 66128 24556 66134 24608
rect 65412 24506 74980 24528
rect 65412 24454 71858 24506
rect 71910 24454 71922 24506
rect 71974 24454 71986 24506
rect 72038 24454 72050 24506
rect 72102 24454 72114 24506
rect 72166 24454 74980 24506
rect 65412 24432 74980 24454
rect 65886 24352 65892 24404
rect 65944 24352 65950 24404
rect 65978 24352 65984 24404
rect 66036 24392 66042 24404
rect 66625 24395 66683 24401
rect 66625 24392 66637 24395
rect 66036 24364 66637 24392
rect 66036 24352 66042 24364
rect 66625 24361 66637 24364
rect 66671 24361 66683 24395
rect 66625 24355 66683 24361
rect 64874 24324 64880 24336
rect 63328 24296 64880 24324
rect 64874 24284 64880 24296
rect 64932 24284 64938 24336
rect 67266 24284 67272 24336
rect 67324 24324 67330 24336
rect 67634 24324 67640 24336
rect 67324 24296 67640 24324
rect 67324 24284 67330 24296
rect 67634 24284 67640 24296
rect 67692 24284 67698 24336
rect 66070 24148 66076 24200
rect 66128 24188 66134 24200
rect 66441 24191 66499 24197
rect 66441 24188 66453 24191
rect 66128 24160 66453 24188
rect 66128 24148 66134 24160
rect 66441 24157 66453 24160
rect 66487 24157 66499 24191
rect 66441 24151 66499 24157
rect 67266 24148 67272 24200
rect 67324 24148 67330 24200
rect 65797 24055 65855 24061
rect 65797 24021 65809 24055
rect 65843 24052 65855 24055
rect 65886 24052 65892 24064
rect 65843 24024 65892 24052
rect 65843 24021 65855 24024
rect 65797 24015 65855 24021
rect 65886 24012 65892 24024
rect 65944 24052 65950 24064
rect 66162 24052 66168 24064
rect 65944 24024 66168 24052
rect 65944 24012 65950 24024
rect 66162 24012 66168 24024
rect 66220 24012 66226 24064
rect 65412 23962 74980 23984
rect 65412 23910 74210 23962
rect 74262 23910 74274 23962
rect 74326 23910 74338 23962
rect 74390 23910 74402 23962
rect 74454 23910 74466 23962
rect 74518 23910 74980 23962
rect 65412 23888 74980 23910
rect 65705 23851 65763 23857
rect 65705 23817 65717 23851
rect 65751 23848 65763 23851
rect 65794 23848 65800 23860
rect 65751 23820 65800 23848
rect 65751 23817 65763 23820
rect 65705 23811 65763 23817
rect 65794 23808 65800 23820
rect 65852 23808 65858 23860
rect 66438 23808 66444 23860
rect 66496 23808 66502 23860
rect 67174 23808 67180 23860
rect 67232 23808 67238 23860
rect 65242 23740 65248 23792
rect 65300 23780 65306 23792
rect 66162 23780 66168 23792
rect 65300 23752 66168 23780
rect 65300 23740 65306 23752
rect 66162 23740 66168 23752
rect 66220 23740 66226 23792
rect 63236 23644 63264 23650
rect 63236 23616 63540 23644
rect 63512 23576 63540 23616
rect 65334 23604 65340 23656
rect 65392 23644 65398 23656
rect 66257 23647 66315 23653
rect 66257 23644 66269 23647
rect 65392 23616 66269 23644
rect 65392 23604 65398 23616
rect 66257 23613 66269 23616
rect 66303 23613 66315 23647
rect 66257 23607 66315 23613
rect 67085 23647 67143 23653
rect 67085 23613 67097 23647
rect 67131 23644 67143 23647
rect 67174 23644 67180 23656
rect 67131 23616 67180 23644
rect 67131 23613 67143 23616
rect 67085 23607 67143 23613
rect 67174 23604 67180 23616
rect 67232 23604 67238 23656
rect 67726 23604 67732 23656
rect 67784 23604 67790 23656
rect 67818 23576 67824 23588
rect 63512 23548 67824 23576
rect 67818 23536 67824 23548
rect 67876 23536 67882 23588
rect 65412 23418 74980 23440
rect 63236 23100 63264 23398
rect 65412 23366 71858 23418
rect 71910 23366 71922 23418
rect 71974 23366 71986 23418
rect 72038 23366 72050 23418
rect 72102 23366 72114 23418
rect 72166 23366 74980 23418
rect 65412 23344 74980 23366
rect 63678 23264 63684 23316
rect 63736 23304 63742 23316
rect 65889 23307 65947 23313
rect 65889 23304 65901 23307
rect 63736 23276 65901 23304
rect 63736 23264 63742 23276
rect 65889 23273 65901 23276
rect 65935 23273 65947 23307
rect 65889 23267 65947 23273
rect 66625 23307 66683 23313
rect 66625 23273 66637 23307
rect 66671 23304 66683 23307
rect 67542 23304 67548 23316
rect 66671 23276 67548 23304
rect 66671 23273 66683 23276
rect 66625 23267 66683 23273
rect 67542 23264 67548 23276
rect 67600 23264 67606 23316
rect 66254 23196 66260 23248
rect 66312 23236 66318 23248
rect 67266 23236 67272 23248
rect 66312 23208 67272 23236
rect 66312 23196 66318 23208
rect 67266 23196 67272 23208
rect 67324 23196 67330 23248
rect 63678 23100 63684 23112
rect 63236 23072 63684 23100
rect 63678 23060 63684 23072
rect 63736 23060 63742 23112
rect 66530 23060 66536 23112
rect 66588 23060 66594 23112
rect 67174 23060 67180 23112
rect 67232 23060 67238 23112
rect 67634 23060 67640 23112
rect 67692 23100 67698 23112
rect 67818 23100 67824 23112
rect 67692 23072 67824 23100
rect 67692 23060 67698 23072
rect 67818 23060 67824 23072
rect 67876 23060 67882 23112
rect 65334 22924 65340 22976
rect 65392 22964 65398 22976
rect 65705 22967 65763 22973
rect 65705 22964 65717 22967
rect 65392 22936 65717 22964
rect 65392 22924 65398 22936
rect 65705 22933 65717 22936
rect 65751 22933 65763 22967
rect 65705 22927 65763 22933
rect 65412 22874 74980 22896
rect 65412 22822 74210 22874
rect 74262 22822 74274 22874
rect 74326 22822 74338 22874
rect 74390 22822 74402 22874
rect 74454 22822 74466 22874
rect 74518 22822 74980 22874
rect 65412 22800 74980 22822
rect 63494 22720 63500 22772
rect 63552 22760 63558 22772
rect 65705 22763 65763 22769
rect 65705 22760 65717 22763
rect 63552 22732 65717 22760
rect 63552 22720 63558 22732
rect 65705 22729 65717 22732
rect 65751 22729 65763 22763
rect 65705 22723 65763 22729
rect 63494 22556 63500 22568
rect 63236 22528 63500 22556
rect 63236 22422 63264 22528
rect 63494 22516 63500 22528
rect 63552 22556 63558 22568
rect 64874 22556 64880 22568
rect 63552 22528 64880 22556
rect 63552 22516 63558 22528
rect 64874 22516 64880 22528
rect 64932 22516 64938 22568
rect 66254 22516 66260 22568
rect 66312 22516 66318 22568
rect 64506 22312 64512 22364
rect 64564 22312 64570 22364
rect 64598 22312 64604 22364
rect 64656 22352 64662 22364
rect 64874 22352 64880 22364
rect 64656 22324 64880 22352
rect 64656 22312 64662 22324
rect 64874 22312 64880 22324
rect 64932 22312 64938 22364
rect 65412 22330 74980 22352
rect 64524 22160 64552 22312
rect 65412 22278 71858 22330
rect 71910 22278 71922 22330
rect 71974 22278 71986 22330
rect 72038 22278 72050 22330
rect 72102 22278 72114 22330
rect 72166 22278 74980 22330
rect 65412 22256 74980 22278
rect 64414 22108 64420 22160
rect 64472 22108 64478 22160
rect 64506 22108 64512 22160
rect 64564 22108 64570 22160
rect 64432 22080 64460 22108
rect 64598 22080 64604 22092
rect 64432 22052 64604 22080
rect 64598 22040 64604 22052
rect 64656 22040 64662 22092
rect 64414 21972 64420 22024
rect 64472 22012 64478 22024
rect 64874 22012 64880 22024
rect 64472 21984 64880 22012
rect 64472 21972 64478 21984
rect 64874 21972 64880 21984
rect 64932 21972 64938 22024
rect 65412 21786 74980 21808
rect 65412 21734 74210 21786
rect 74262 21734 74274 21786
rect 74326 21734 74338 21786
rect 74390 21734 74402 21786
rect 74454 21734 74466 21786
rect 74518 21734 74980 21786
rect 65412 21712 74980 21734
rect 63328 21400 63356 21470
rect 70210 21400 70216 21412
rect 63328 21372 70216 21400
rect 70210 21360 70216 21372
rect 70268 21360 70274 21412
rect 63494 21292 63500 21344
rect 63552 21332 63558 21344
rect 63552 21304 63632 21332
rect 63552 21292 63558 21304
rect 63494 21232 63500 21244
rect 63342 21204 63500 21232
rect 63494 21192 63500 21204
rect 63552 21192 63558 21244
rect 63604 20720 63632 21304
rect 65412 21242 74980 21264
rect 65412 21190 71858 21242
rect 71910 21190 71922 21242
rect 71974 21190 71986 21242
rect 72038 21190 72050 21242
rect 72102 21190 72114 21242
rect 72166 21190 74980 21242
rect 65412 21168 74980 21190
rect 63328 20692 63632 20720
rect 65412 20698 74980 20720
rect 63328 19428 63356 20692
rect 65412 20646 74210 20698
rect 74262 20646 74274 20698
rect 74326 20646 74338 20698
rect 74390 20646 74402 20698
rect 74454 20646 74466 20698
rect 74518 20646 74980 20698
rect 65412 20624 74980 20646
rect 65412 20154 74980 20176
rect 65412 20102 71858 20154
rect 71910 20102 71922 20154
rect 71974 20102 71986 20154
rect 72038 20102 72050 20154
rect 72102 20102 72114 20154
rect 72166 20102 74980 20154
rect 65412 20080 74980 20102
rect 65412 19610 74980 19632
rect 65412 19558 74210 19610
rect 74262 19558 74274 19610
rect 74326 19558 74338 19610
rect 74390 19558 74402 19610
rect 74454 19558 74466 19610
rect 74518 19558 74980 19610
rect 65412 19536 74980 19558
rect 63328 19400 63632 19428
rect 63604 19292 63632 19400
rect 64874 19292 64880 19304
rect 63328 19156 63356 19290
rect 63604 19264 64880 19292
rect 64874 19252 64880 19264
rect 64932 19252 64938 19304
rect 66254 19156 66260 19168
rect 63328 19128 66260 19156
rect 66254 19116 66260 19128
rect 66312 19116 66318 19168
rect 65412 19066 74980 19088
rect 63328 18884 63356 19038
rect 65412 19014 71858 19066
rect 71910 19014 71922 19066
rect 71974 19014 71986 19066
rect 72038 19014 72050 19066
rect 72102 19014 72114 19066
rect 72166 19014 74980 19066
rect 65412 18992 74980 19014
rect 67818 18952 67824 18964
rect 67606 18924 67824 18952
rect 67606 18884 67634 18924
rect 67818 18912 67824 18924
rect 67876 18912 67882 18964
rect 63328 18856 67634 18884
rect 65412 18522 74980 18544
rect 65412 18470 74210 18522
rect 74262 18470 74274 18522
rect 74326 18470 74338 18522
rect 74390 18470 74402 18522
rect 74454 18470 74466 18522
rect 74518 18470 74980 18522
rect 65412 18448 74980 18470
rect 63678 18068 63684 18080
rect 63328 18040 63684 18068
rect 63678 18028 63684 18040
rect 63736 18068 63742 18080
rect 64874 18068 64880 18080
rect 63736 18040 64880 18068
rect 63736 18028 63742 18040
rect 64874 18028 64880 18040
rect 64932 18028 64938 18080
rect 65412 17978 74980 18000
rect 65412 17926 71858 17978
rect 71910 17926 71922 17978
rect 71974 17926 71986 17978
rect 72038 17926 72050 17978
rect 72102 17926 72114 17978
rect 72166 17926 74980 17978
rect 65412 17904 74980 17926
rect 64598 17552 64604 17604
rect 64656 17592 64662 17604
rect 65058 17592 65064 17604
rect 64656 17564 65064 17592
rect 64656 17552 64662 17564
rect 65058 17552 65064 17564
rect 65116 17552 65122 17604
rect 64138 17416 64144 17468
rect 64196 17456 64202 17468
rect 64598 17456 64604 17468
rect 64196 17428 64604 17456
rect 64196 17416 64202 17428
rect 64598 17416 64604 17428
rect 64656 17416 64662 17468
rect 65412 17434 74980 17456
rect 65412 17382 74210 17434
rect 74262 17382 74274 17434
rect 74326 17382 74338 17434
rect 74390 17382 74402 17434
rect 74454 17382 74466 17434
rect 74518 17382 74980 17434
rect 65412 17360 74980 17382
rect 66530 17212 66536 17264
rect 66588 17252 66594 17264
rect 66806 17252 66812 17264
rect 66588 17224 66812 17252
rect 66588 17212 66594 17224
rect 66806 17212 66812 17224
rect 66864 17212 66870 17264
rect 63328 16980 63356 17110
rect 63328 16952 63448 16980
rect 63328 16640 63356 16858
rect 63420 16776 63448 16952
rect 65412 16890 74980 16912
rect 65412 16838 71858 16890
rect 71910 16838 71922 16890
rect 71974 16838 71986 16890
rect 72038 16838 72050 16890
rect 72102 16838 72114 16890
rect 72166 16838 74980 16890
rect 65412 16816 74980 16838
rect 65886 16776 65892 16788
rect 63420 16748 65892 16776
rect 65886 16736 65892 16748
rect 65944 16736 65950 16788
rect 65978 16640 65984 16652
rect 63328 16612 65984 16640
rect 65978 16600 65984 16612
rect 66036 16600 66042 16652
rect 65412 16346 74980 16368
rect 65412 16294 74210 16346
rect 74262 16294 74274 16346
rect 74326 16294 74338 16346
rect 74390 16294 74402 16346
rect 74454 16294 74466 16346
rect 74518 16294 74980 16346
rect 65412 16272 74980 16294
rect 63328 15620 63356 15882
rect 65412 15802 74980 15824
rect 65412 15750 71858 15802
rect 71910 15750 71922 15802
rect 71974 15750 71986 15802
rect 72038 15750 72050 15802
rect 72102 15750 72114 15802
rect 72166 15750 74980 15802
rect 65412 15728 74980 15750
rect 63586 15620 63592 15632
rect 63328 15592 63592 15620
rect 63586 15580 63592 15592
rect 63644 15580 63650 15632
rect 65412 15258 74980 15280
rect 65412 15206 74210 15258
rect 74262 15206 74274 15258
rect 74326 15206 74338 15258
rect 74390 15206 74402 15258
rect 74454 15206 74466 15258
rect 74518 15206 74980 15258
rect 65412 15184 74980 15206
rect 63328 14804 63356 14930
rect 66806 14804 66812 14816
rect 63328 14776 66812 14804
rect 66806 14764 66812 14776
rect 66864 14764 66870 14816
rect 65412 14714 74980 14736
rect 63328 14396 63356 14678
rect 65412 14662 71858 14714
rect 71910 14662 71922 14714
rect 71974 14662 71986 14714
rect 72038 14662 72050 14714
rect 72102 14662 72114 14714
rect 72166 14662 74980 14714
rect 65412 14640 74980 14662
rect 65242 14396 65248 14408
rect 63328 14368 65248 14396
rect 65242 14356 65248 14368
rect 65300 14356 65306 14408
rect 65412 14170 74980 14192
rect 65412 14118 74210 14170
rect 74262 14118 74274 14170
rect 74326 14118 74338 14170
rect 74390 14118 74402 14170
rect 74454 14118 74466 14170
rect 74518 14118 74980 14170
rect 65412 14096 74980 14118
rect 63586 13716 63592 13728
rect 63342 13688 63592 13716
rect 63586 13676 63592 13688
rect 63644 13676 63650 13728
rect 65412 13626 74980 13648
rect 65412 13574 71858 13626
rect 71910 13574 71922 13626
rect 71974 13574 71986 13626
rect 72038 13574 72050 13626
rect 72102 13574 72114 13626
rect 72166 13574 74980 13626
rect 65412 13552 74980 13574
rect 65412 13082 74980 13104
rect 65412 13030 74210 13082
rect 74262 13030 74274 13082
rect 74326 13030 74338 13082
rect 74390 13030 74402 13082
rect 74454 13030 74466 13082
rect 74518 13030 74980 13082
rect 65412 13008 74980 13030
rect 63328 12628 63356 12750
rect 66070 12628 66076 12640
rect 63328 12600 66076 12628
rect 66070 12588 66076 12600
rect 66128 12588 66134 12640
rect 65412 12538 74980 12560
rect 63328 12492 63356 12498
rect 64874 12492 64880 12504
rect 63328 12464 64880 12492
rect 64874 12452 64880 12464
rect 64932 12452 64938 12504
rect 65412 12486 71858 12538
rect 71910 12486 71922 12538
rect 71974 12486 71986 12538
rect 72038 12486 72050 12538
rect 72102 12486 72114 12538
rect 72166 12486 74980 12538
rect 65412 12464 74980 12486
rect 63678 12384 63684 12436
rect 63736 12424 63742 12436
rect 65058 12424 65064 12436
rect 63736 12396 65064 12424
rect 63736 12384 63742 12396
rect 65058 12384 65064 12396
rect 65116 12384 65122 12436
rect 63954 11976 63960 12028
rect 64012 12016 64018 12028
rect 64782 12016 64788 12028
rect 64012 11988 64788 12016
rect 64012 11976 64018 11988
rect 64782 11976 64788 11988
rect 64840 11976 64846 12028
rect 65412 11994 74980 12016
rect 65412 11942 74210 11994
rect 74262 11942 74274 11994
rect 74326 11942 74338 11994
rect 74390 11942 74402 11994
rect 74454 11942 74466 11994
rect 74518 11942 74980 11994
rect 65412 11920 74980 11942
rect 64598 11840 64604 11892
rect 64656 11880 64662 11892
rect 64782 11880 64788 11892
rect 64656 11852 64788 11880
rect 64656 11840 64662 11852
rect 64782 11840 64788 11852
rect 64840 11840 64846 11892
rect 65058 11840 65064 11892
rect 65116 11880 65122 11892
rect 65334 11880 65340 11892
rect 65116 11852 65340 11880
rect 65116 11840 65122 11852
rect 65334 11840 65340 11852
rect 65392 11840 65398 11892
rect 63586 11540 63592 11552
rect 63328 11512 63592 11540
rect 63586 11500 63592 11512
rect 63644 11500 63650 11552
rect 65412 11450 74980 11472
rect 65412 11398 71858 11450
rect 71910 11398 71922 11450
rect 71974 11398 71986 11450
rect 72038 11398 72050 11450
rect 72102 11398 72114 11450
rect 72166 11398 74980 11450
rect 65412 11376 74980 11398
rect 65412 10906 74980 10928
rect 65412 10854 74210 10906
rect 74262 10854 74274 10906
rect 74326 10854 74338 10906
rect 74390 10854 74402 10906
rect 74454 10854 74466 10906
rect 74518 10854 74980 10906
rect 65412 10832 74980 10854
rect 63328 10696 64184 10724
rect 63328 10588 63356 10696
rect 63236 10560 63356 10588
rect 63328 10248 63356 10318
rect 63586 10292 63592 10344
rect 63644 10292 63650 10344
rect 63604 10248 63632 10292
rect 63328 10220 63632 10248
rect 64156 10248 64184 10696
rect 66530 10684 66536 10736
rect 66588 10724 66594 10736
rect 67174 10724 67180 10736
rect 66588 10696 67180 10724
rect 66588 10684 66594 10696
rect 67174 10684 67180 10696
rect 67232 10684 67238 10736
rect 66806 10548 66812 10600
rect 66864 10588 66870 10600
rect 67174 10588 67180 10600
rect 66864 10560 67180 10588
rect 66864 10548 66870 10560
rect 67174 10548 67180 10560
rect 67232 10548 67238 10600
rect 65412 10362 74980 10384
rect 65412 10310 71858 10362
rect 71910 10310 71922 10362
rect 71974 10310 71986 10362
rect 72038 10310 72050 10362
rect 72102 10310 72114 10362
rect 72166 10310 74980 10362
rect 65412 10288 74980 10310
rect 66806 10248 66812 10260
rect 64156 10220 66812 10248
rect 66806 10208 66812 10220
rect 66864 10208 66870 10260
rect 63494 10004 63500 10056
rect 63552 10044 63558 10056
rect 63552 10016 63632 10044
rect 63552 10004 63558 10016
rect 63604 9704 63632 10016
rect 65412 9818 74980 9840
rect 65412 9766 74210 9818
rect 74262 9766 74274 9818
rect 74326 9766 74338 9818
rect 74390 9766 74402 9818
rect 74454 9766 74466 9818
rect 74518 9766 74980 9818
rect 65412 9744 74980 9766
rect 63328 9676 63632 9704
rect 63328 9342 63356 9676
rect 65412 9274 74980 9296
rect 65412 9222 71858 9274
rect 71910 9222 71922 9274
rect 71974 9222 71986 9274
rect 72038 9222 72050 9274
rect 72102 9222 72114 9274
rect 72166 9222 74980 9274
rect 65412 9200 74980 9222
rect 65426 9120 65432 9172
rect 65484 9160 65490 9172
rect 65484 9132 66116 9160
rect 65484 9120 65490 9132
rect 65426 8984 65432 9036
rect 65484 9024 65490 9036
rect 65978 9024 65984 9036
rect 65484 8996 65984 9024
rect 65484 8984 65490 8996
rect 65978 8984 65984 8996
rect 66036 8984 66042 9036
rect 66088 8832 66116 9132
rect 66070 8780 66076 8832
rect 66128 8780 66134 8832
rect 65412 8730 74980 8752
rect 65412 8678 74210 8730
rect 74262 8678 74274 8730
rect 74326 8678 74338 8730
rect 74390 8678 74402 8730
rect 74454 8678 74466 8730
rect 74518 8678 74980 8730
rect 65412 8656 74980 8678
rect 66438 8276 66444 8288
rect 63052 8248 66444 8276
rect 63052 7936 63080 8248
rect 66438 8236 66444 8248
rect 66496 8236 66502 8288
rect 65412 8186 74980 8208
rect 65412 8134 71858 8186
rect 71910 8134 71922 8186
rect 71974 8134 71986 8186
rect 72038 8134 72050 8186
rect 72102 8134 72114 8186
rect 72166 8134 74980 8186
rect 65412 8112 74980 8134
rect 66438 8032 66444 8084
rect 66496 8072 66502 8084
rect 66898 8072 66904 8084
rect 66496 8044 66904 8072
rect 66496 8032 66502 8044
rect 66898 8032 66904 8044
rect 66956 8032 66962 8084
rect 67726 8032 67732 8084
rect 67784 8032 67790 8084
rect 64230 7936 64236 7948
rect 50724 7908 60734 7936
rect 50724 7880 50752 7908
rect 50706 7828 50712 7880
rect 50764 7828 50770 7880
rect 60706 7800 60734 7908
rect 62960 7908 63080 7936
rect 63144 7908 64236 7936
rect 62482 7828 62488 7880
rect 62540 7868 62546 7880
rect 62960 7868 62988 7908
rect 62540 7840 62988 7868
rect 62540 7828 62546 7840
rect 63144 7800 63172 7908
rect 64230 7896 64236 7908
rect 64288 7896 64294 7948
rect 63218 7828 63224 7880
rect 63276 7868 63282 7880
rect 67744 7868 67772 8032
rect 67910 7896 67916 7948
rect 67968 7936 67974 7948
rect 68646 7936 68652 7948
rect 67968 7908 68652 7936
rect 67968 7896 67974 7908
rect 68646 7896 68652 7908
rect 68704 7896 68710 7948
rect 63276 7840 67772 7868
rect 63276 7828 63282 7840
rect 60706 7772 63172 7800
rect 63402 7760 63408 7812
rect 63460 7800 63466 7812
rect 66346 7800 66352 7812
rect 63460 7772 66352 7800
rect 63460 7760 63466 7772
rect 66346 7760 66352 7772
rect 66404 7760 66410 7812
rect 66438 7760 66444 7812
rect 66496 7760 66502 7812
rect 66530 7760 66536 7812
rect 66588 7800 66594 7812
rect 66990 7800 66996 7812
rect 66588 7772 66996 7800
rect 66588 7760 66594 7772
rect 66990 7760 66996 7772
rect 67048 7760 67054 7812
rect 35986 7692 35992 7744
rect 36044 7732 36050 7744
rect 64046 7732 64052 7744
rect 36044 7704 64052 7732
rect 36044 7692 36050 7704
rect 64046 7692 64052 7704
rect 64104 7692 64110 7744
rect 66456 7732 66484 7760
rect 64248 7704 66484 7732
rect 36078 7624 36084 7676
rect 36136 7664 36142 7676
rect 64138 7664 64144 7676
rect 36136 7636 64144 7664
rect 36136 7624 36142 7636
rect 64138 7624 64144 7636
rect 64196 7624 64202 7676
rect 32950 7556 32956 7608
rect 33008 7596 33014 7608
rect 63678 7596 63684 7608
rect 33008 7568 63684 7596
rect 33008 7556 33014 7568
rect 63678 7556 63684 7568
rect 63736 7556 63742 7608
rect 58986 7488 58992 7540
rect 59044 7528 59050 7540
rect 64248 7528 64276 7704
rect 65412 7642 74980 7664
rect 65412 7590 74210 7642
rect 74262 7590 74274 7642
rect 74326 7590 74338 7642
rect 74390 7590 74402 7642
rect 74454 7590 74466 7642
rect 74518 7590 74980 7642
rect 65412 7568 74980 7590
rect 59044 7500 64276 7528
rect 59044 7488 59050 7500
rect 64782 7488 64788 7540
rect 64840 7528 64846 7540
rect 65705 7531 65763 7537
rect 65705 7528 65717 7531
rect 64840 7500 65717 7528
rect 64840 7488 64846 7500
rect 65705 7497 65717 7500
rect 65751 7497 65763 7531
rect 65705 7491 65763 7497
rect 69198 7488 69204 7540
rect 69256 7488 69262 7540
rect 59998 7352 60004 7404
rect 60056 7392 60062 7404
rect 65794 7392 65800 7404
rect 60056 7364 65800 7392
rect 60056 7352 60062 7364
rect 65794 7352 65800 7364
rect 65852 7352 65858 7404
rect 66530 7352 66536 7404
rect 66588 7392 66594 7404
rect 67082 7392 67088 7404
rect 66588 7364 67088 7392
rect 66588 7352 66594 7364
rect 67082 7352 67088 7364
rect 67140 7352 67146 7404
rect 58894 7284 58900 7336
rect 58952 7324 58958 7336
rect 65426 7324 65432 7336
rect 58952 7296 65432 7324
rect 58952 7284 58958 7296
rect 65426 7284 65432 7296
rect 65484 7284 65490 7336
rect 59078 7216 59084 7268
rect 59136 7256 59142 7268
rect 65978 7256 65984 7268
rect 59136 7228 65984 7256
rect 59136 7216 59142 7228
rect 65978 7216 65984 7228
rect 66036 7216 66042 7268
rect 59538 7148 59544 7200
rect 59596 7188 59602 7200
rect 66806 7188 66812 7200
rect 59596 7160 66812 7188
rect 59596 7148 59602 7160
rect 66806 7148 66812 7160
rect 66864 7148 66870 7200
rect 59262 7080 59268 7132
rect 59320 7120 59326 7132
rect 65150 7120 65156 7132
rect 59320 7092 65156 7120
rect 59320 7080 59326 7092
rect 65150 7080 65156 7092
rect 65208 7080 65214 7132
rect 65412 7098 74980 7120
rect 59722 7012 59728 7064
rect 59780 7052 59786 7064
rect 63954 7052 63960 7064
rect 59780 7024 63960 7052
rect 59780 7012 59786 7024
rect 63954 7012 63960 7024
rect 64012 7012 64018 7064
rect 65412 7046 71858 7098
rect 71910 7046 71922 7098
rect 71974 7046 71986 7098
rect 72038 7046 72050 7098
rect 72102 7046 72114 7098
rect 72166 7046 74980 7098
rect 65412 7024 74980 7046
rect 59354 6944 59360 6996
rect 59412 6984 59418 6996
rect 65334 6984 65340 6996
rect 59412 6956 65340 6984
rect 59412 6944 59418 6956
rect 65334 6944 65340 6956
rect 65392 6944 65398 6996
rect 66530 6944 66536 6996
rect 66588 6944 66594 6996
rect 69198 6944 69204 6996
rect 69256 6944 69262 6996
rect 61194 6876 61200 6928
rect 61252 6916 61258 6928
rect 63494 6916 63500 6928
rect 61252 6888 63500 6916
rect 61252 6876 61258 6888
rect 63494 6876 63500 6888
rect 63552 6876 63558 6928
rect 48130 6808 48136 6860
rect 48188 6848 48194 6860
rect 48188 6820 64552 6848
rect 48188 6808 48194 6820
rect 36630 6740 36636 6792
rect 36688 6780 36694 6792
rect 64230 6780 64236 6792
rect 36688 6752 64236 6780
rect 36688 6740 36694 6752
rect 64230 6740 64236 6752
rect 64288 6740 64294 6792
rect 64524 6780 64552 6820
rect 64598 6808 64604 6860
rect 64656 6848 64662 6860
rect 67450 6848 67456 6860
rect 64656 6820 67456 6848
rect 64656 6808 64662 6820
rect 67450 6808 67456 6820
rect 67508 6808 67514 6860
rect 69290 6780 69296 6792
rect 64524 6752 69296 6780
rect 69290 6740 69296 6752
rect 69348 6740 69354 6792
rect 35158 6672 35164 6724
rect 35216 6712 35222 6724
rect 62850 6712 62856 6724
rect 35216 6684 62856 6712
rect 35216 6672 35222 6684
rect 62850 6672 62856 6684
rect 62908 6672 62914 6724
rect 51442 6604 51448 6656
rect 51500 6644 51506 6656
rect 68462 6644 68468 6656
rect 51500 6616 68468 6644
rect 51500 6604 51506 6616
rect 68462 6604 68468 6616
rect 68520 6604 68526 6656
rect 33686 6536 33692 6588
rect 33744 6576 33750 6588
rect 64506 6576 64512 6588
rect 33744 6548 64512 6576
rect 33744 6536 33750 6548
rect 64506 6536 64512 6548
rect 64564 6536 64570 6588
rect 65412 6554 74980 6576
rect 30466 6468 30472 6520
rect 30524 6508 30530 6520
rect 30524 6480 64552 6508
rect 65412 6502 74210 6554
rect 74262 6502 74274 6554
rect 74326 6502 74338 6554
rect 74390 6502 74402 6554
rect 74454 6502 74466 6554
rect 74518 6502 74980 6554
rect 65412 6480 74980 6502
rect 30524 6468 30530 6480
rect 30282 6400 30288 6452
rect 30340 6440 30346 6452
rect 30340 6412 48314 6440
rect 30340 6400 30346 6412
rect 31018 6332 31024 6384
rect 31076 6372 31082 6384
rect 48286 6372 48314 6412
rect 52270 6400 52276 6452
rect 52328 6440 52334 6452
rect 64414 6440 64420 6452
rect 52328 6412 64420 6440
rect 52328 6400 52334 6412
rect 64414 6400 64420 6412
rect 64472 6400 64478 6452
rect 64524 6440 64552 6480
rect 65886 6440 65892 6452
rect 64524 6412 65892 6440
rect 65886 6400 65892 6412
rect 65944 6400 65950 6452
rect 66530 6400 66536 6452
rect 66588 6400 66594 6452
rect 69198 6400 69204 6452
rect 69256 6400 69262 6452
rect 31076 6344 41414 6372
rect 48286 6344 52408 6372
rect 31076 6332 31082 6344
rect 41386 6236 41414 6344
rect 52380 6304 52408 6344
rect 53098 6332 53104 6384
rect 53156 6372 53162 6384
rect 62758 6372 62764 6384
rect 53156 6344 62764 6372
rect 53156 6332 53162 6344
rect 62758 6332 62764 6344
rect 62816 6332 62822 6384
rect 62850 6332 62856 6384
rect 62908 6372 62914 6384
rect 69382 6372 69388 6384
rect 62908 6344 69388 6372
rect 62908 6332 62914 6344
rect 69382 6332 69388 6344
rect 69440 6332 69446 6384
rect 67174 6304 67180 6316
rect 52380 6276 67180 6304
rect 67174 6264 67180 6276
rect 67232 6264 67238 6316
rect 53098 6236 53104 6248
rect 41386 6208 53104 6236
rect 53098 6196 53104 6208
rect 53156 6196 53162 6248
rect 56594 6196 56600 6248
rect 56652 6236 56658 6248
rect 64874 6236 64880 6248
rect 56652 6208 64880 6236
rect 56652 6196 56658 6208
rect 64874 6196 64880 6208
rect 64932 6196 64938 6248
rect 47302 6128 47308 6180
rect 47360 6168 47366 6180
rect 65518 6168 65524 6180
rect 47360 6140 65524 6168
rect 47360 6128 47366 6140
rect 65518 6128 65524 6140
rect 65576 6128 65582 6180
rect 65886 6128 65892 6180
rect 65944 6168 65950 6180
rect 69014 6168 69020 6180
rect 65944 6140 69020 6168
rect 65944 6128 65950 6140
rect 69014 6128 69020 6140
rect 69072 6128 69078 6180
rect 53282 6060 53288 6112
rect 53340 6100 53346 6112
rect 61470 6100 61476 6112
rect 53340 6072 61476 6100
rect 53340 6060 53346 6072
rect 61470 6060 61476 6072
rect 61528 6060 61534 6112
rect 62758 6060 62764 6112
rect 62816 6100 62822 6112
rect 64046 6100 64052 6112
rect 62816 6072 64052 6100
rect 62816 6060 62822 6072
rect 64046 6060 64052 6072
rect 64104 6060 64110 6112
rect 64230 6060 64236 6112
rect 64288 6100 64294 6112
rect 69566 6100 69572 6112
rect 64288 6072 69572 6100
rect 64288 6060 64294 6072
rect 69566 6060 69572 6072
rect 69624 6060 69630 6112
rect 1012 6010 74980 6032
rect 1012 5958 71858 6010
rect 71910 5958 71922 6010
rect 71974 5958 71986 6010
rect 72038 5958 72050 6010
rect 72102 5958 72114 6010
rect 72166 5958 74980 6010
rect 1012 5936 74980 5958
rect 50706 5856 50712 5908
rect 50764 5856 50770 5908
rect 51442 5856 51448 5908
rect 51500 5856 51506 5908
rect 52181 5899 52239 5905
rect 52181 5865 52193 5899
rect 52227 5896 52239 5899
rect 52270 5896 52276 5908
rect 52227 5868 52276 5896
rect 52227 5865 52239 5868
rect 52181 5859 52239 5865
rect 52270 5856 52276 5868
rect 52328 5856 52334 5908
rect 53282 5856 53288 5908
rect 53340 5856 53346 5908
rect 55861 5899 55919 5905
rect 55861 5865 55873 5899
rect 55907 5896 55919 5899
rect 55907 5868 58296 5896
rect 55907 5865 55919 5868
rect 55861 5859 55919 5865
rect 42702 5788 42708 5840
rect 42760 5788 42766 5840
rect 44726 5788 44732 5840
rect 44784 5788 44790 5840
rect 54757 5831 54815 5837
rect 54757 5797 54769 5831
rect 54803 5828 54815 5831
rect 58268 5828 58296 5868
rect 59170 5856 59176 5908
rect 59228 5896 59234 5908
rect 59357 5899 59415 5905
rect 59357 5896 59369 5899
rect 59228 5868 59369 5896
rect 59228 5856 59234 5868
rect 59357 5865 59369 5868
rect 59403 5896 59415 5899
rect 59541 5899 59599 5905
rect 59541 5896 59553 5899
rect 59403 5868 59553 5896
rect 59403 5865 59415 5868
rect 59357 5859 59415 5865
rect 59541 5865 59553 5868
rect 59587 5896 59599 5899
rect 59722 5896 59728 5908
rect 59587 5868 59728 5896
rect 59587 5865 59599 5868
rect 59541 5859 59599 5865
rect 59722 5856 59728 5868
rect 59780 5856 59786 5908
rect 60645 5899 60703 5905
rect 60645 5865 60657 5899
rect 60691 5896 60703 5899
rect 60734 5896 60740 5908
rect 60691 5868 60740 5896
rect 60691 5865 60703 5868
rect 60645 5859 60703 5865
rect 60734 5856 60740 5868
rect 60792 5896 60798 5908
rect 60829 5899 60887 5905
rect 60829 5896 60841 5899
rect 60792 5868 60841 5896
rect 60792 5856 60798 5868
rect 60829 5865 60841 5868
rect 60875 5896 60887 5899
rect 61013 5899 61071 5905
rect 61013 5896 61025 5899
rect 60875 5868 61025 5896
rect 60875 5865 60887 5868
rect 60829 5859 60887 5865
rect 61013 5865 61025 5868
rect 61059 5896 61071 5899
rect 61194 5896 61200 5908
rect 61059 5868 61200 5896
rect 61059 5865 61071 5868
rect 61013 5859 61071 5865
rect 61194 5856 61200 5868
rect 61252 5856 61258 5908
rect 61286 5856 61292 5908
rect 61344 5896 61350 5908
rect 63494 5896 63500 5908
rect 61344 5868 63500 5896
rect 61344 5856 61350 5868
rect 63494 5856 63500 5868
rect 63552 5856 63558 5908
rect 63586 5856 63592 5908
rect 63644 5896 63650 5908
rect 63773 5899 63831 5905
rect 63773 5896 63785 5899
rect 63644 5868 63785 5896
rect 63644 5856 63650 5868
rect 63773 5865 63785 5868
rect 63819 5896 63831 5899
rect 63957 5899 64015 5905
rect 63957 5896 63969 5899
rect 63819 5868 63969 5896
rect 63819 5865 63831 5868
rect 63773 5859 63831 5865
rect 63957 5865 63969 5868
rect 64003 5896 64015 5899
rect 64782 5896 64788 5908
rect 64003 5868 64788 5896
rect 64003 5865 64015 5868
rect 63957 5859 64015 5865
rect 64782 5856 64788 5868
rect 64840 5856 64846 5908
rect 66530 5856 66536 5908
rect 66588 5856 66594 5908
rect 69198 5856 69204 5908
rect 69256 5856 69262 5908
rect 65242 5828 65248 5840
rect 54803 5800 57744 5828
rect 58268 5800 65248 5828
rect 54803 5797 54815 5800
rect 54757 5791 54815 5797
rect 49605 5763 49663 5769
rect 49605 5729 49617 5763
rect 49651 5760 49663 5763
rect 49651 5732 56824 5760
rect 49651 5729 49663 5732
rect 49605 5723 49663 5729
rect 31110 5652 31116 5704
rect 31168 5692 31174 5704
rect 34790 5692 34796 5704
rect 31168 5664 34796 5692
rect 31168 5652 31174 5664
rect 34790 5652 34796 5664
rect 34848 5692 34854 5704
rect 35894 5692 35900 5704
rect 34848 5664 35900 5692
rect 34848 5652 34854 5664
rect 35894 5652 35900 5664
rect 35952 5652 35958 5704
rect 41506 5652 41512 5704
rect 41564 5692 41570 5704
rect 42518 5692 42524 5704
rect 41564 5664 42524 5692
rect 41564 5652 41570 5664
rect 42518 5652 42524 5664
rect 42576 5652 42582 5704
rect 44085 5695 44143 5701
rect 44085 5661 44097 5695
rect 44131 5661 44143 5695
rect 44085 5655 44143 5661
rect 33226 5584 33232 5636
rect 33284 5624 33290 5636
rect 43901 5627 43959 5633
rect 43901 5624 43913 5627
rect 33284 5596 43913 5624
rect 33284 5584 33290 5596
rect 43901 5593 43913 5596
rect 43947 5624 43959 5627
rect 44100 5624 44128 5655
rect 45554 5652 45560 5704
rect 45612 5652 45618 5704
rect 48961 5695 49019 5701
rect 48961 5692 48973 5695
rect 48792 5664 48973 5692
rect 43947 5596 44128 5624
rect 43947 5593 43959 5596
rect 43901 5587 43959 5593
rect 29822 5516 29828 5568
rect 29880 5556 29886 5568
rect 36170 5556 36176 5568
rect 29880 5528 36176 5556
rect 29880 5516 29886 5528
rect 36170 5516 36176 5528
rect 36228 5516 36234 5568
rect 47210 5516 47216 5568
rect 47268 5556 47274 5568
rect 48792 5565 48820 5664
rect 48961 5661 48973 5664
rect 49007 5661 49019 5695
rect 48961 5655 49019 5661
rect 49050 5652 49056 5704
rect 49108 5692 49114 5704
rect 50065 5695 50123 5701
rect 50065 5692 50077 5695
rect 49108 5664 50077 5692
rect 49108 5652 49114 5664
rect 50065 5661 50077 5664
rect 50111 5661 50123 5695
rect 50065 5655 50123 5661
rect 50798 5652 50804 5704
rect 50856 5652 50862 5704
rect 51258 5652 51264 5704
rect 51316 5692 51322 5704
rect 51537 5695 51595 5701
rect 51537 5692 51549 5695
rect 51316 5664 51549 5692
rect 51316 5652 51322 5664
rect 51537 5661 51549 5664
rect 51583 5661 51595 5695
rect 51537 5655 51595 5661
rect 51718 5652 51724 5704
rect 51776 5692 51782 5704
rect 52641 5695 52699 5701
rect 52641 5692 52653 5695
rect 51776 5664 52653 5692
rect 51776 5652 51782 5664
rect 52641 5661 52653 5664
rect 52687 5661 52699 5695
rect 52641 5655 52699 5661
rect 52730 5652 52736 5704
rect 52788 5692 52794 5704
rect 53377 5695 53435 5701
rect 53377 5692 53389 5695
rect 52788 5664 53389 5692
rect 52788 5652 52794 5664
rect 53377 5661 53389 5664
rect 53423 5661 53435 5695
rect 54113 5695 54171 5701
rect 54113 5692 54125 5695
rect 53377 5655 53435 5661
rect 53484 5664 54125 5692
rect 51166 5584 51172 5636
rect 51224 5624 51230 5636
rect 53484 5624 53512 5664
rect 54113 5661 54125 5664
rect 54159 5661 54171 5695
rect 54113 5655 54171 5661
rect 55214 5652 55220 5704
rect 55272 5652 55278 5704
rect 55950 5652 55956 5704
rect 56008 5652 56014 5704
rect 56594 5652 56600 5704
rect 56652 5652 56658 5704
rect 56686 5652 56692 5704
rect 56744 5652 56750 5704
rect 56796 5692 56824 5732
rect 57330 5720 57336 5772
rect 57388 5720 57394 5772
rect 57716 5760 57744 5800
rect 65242 5788 65248 5800
rect 65300 5788 65306 5840
rect 65794 5788 65800 5840
rect 65852 5828 65858 5840
rect 66162 5828 66168 5840
rect 65852 5800 66168 5828
rect 65852 5788 65858 5800
rect 66162 5788 66168 5800
rect 66220 5788 66226 5840
rect 60826 5760 60832 5772
rect 57716 5732 60832 5760
rect 60826 5720 60832 5732
rect 60884 5720 60890 5772
rect 64046 5720 64052 5772
rect 64104 5760 64110 5772
rect 70210 5760 70216 5772
rect 64104 5732 70216 5760
rect 64104 5720 64110 5732
rect 70210 5720 70216 5732
rect 70268 5720 70274 5772
rect 64690 5692 64696 5704
rect 56796 5664 64696 5692
rect 64690 5652 64696 5664
rect 64748 5652 64754 5704
rect 64782 5652 64788 5704
rect 64840 5692 64846 5704
rect 66990 5692 66996 5704
rect 64840 5664 66996 5692
rect 64840 5652 64846 5664
rect 66990 5652 66996 5664
rect 67048 5652 67054 5704
rect 51224 5596 53512 5624
rect 54021 5627 54079 5633
rect 51224 5584 51230 5596
rect 54021 5593 54033 5627
rect 54067 5624 54079 5627
rect 62850 5624 62856 5636
rect 54067 5596 62856 5624
rect 54067 5593 54079 5596
rect 54021 5587 54079 5593
rect 62850 5584 62856 5596
rect 62908 5584 62914 5636
rect 65886 5624 65892 5636
rect 62960 5596 65892 5624
rect 48777 5559 48835 5565
rect 48777 5556 48789 5559
rect 47268 5528 48789 5556
rect 47268 5516 47274 5528
rect 48777 5525 48789 5528
rect 48823 5525 48835 5559
rect 48777 5519 48835 5525
rect 62117 5559 62175 5565
rect 62117 5525 62129 5559
rect 62163 5556 62175 5559
rect 62298 5556 62304 5568
rect 62163 5528 62304 5556
rect 62163 5525 62175 5528
rect 62117 5519 62175 5525
rect 62298 5516 62304 5528
rect 62356 5556 62362 5568
rect 62485 5559 62543 5565
rect 62485 5556 62497 5559
rect 62356 5528 62497 5556
rect 62356 5516 62362 5528
rect 62485 5525 62497 5528
rect 62531 5556 62543 5559
rect 62669 5559 62727 5565
rect 62669 5556 62681 5559
rect 62531 5528 62681 5556
rect 62531 5525 62543 5528
rect 62485 5519 62543 5525
rect 62669 5525 62681 5528
rect 62715 5556 62727 5559
rect 62960 5556 62988 5596
rect 65886 5584 65892 5596
rect 65944 5584 65950 5636
rect 66162 5584 66168 5636
rect 66220 5624 66226 5636
rect 67542 5624 67548 5636
rect 66220 5596 67548 5624
rect 66220 5584 66226 5596
rect 67542 5584 67548 5596
rect 67600 5584 67606 5636
rect 62715 5528 62988 5556
rect 62715 5525 62727 5528
rect 62669 5519 62727 5525
rect 63494 5516 63500 5568
rect 63552 5556 63558 5568
rect 67726 5556 67732 5568
rect 63552 5528 67732 5556
rect 63552 5516 63558 5528
rect 67726 5516 67732 5528
rect 67784 5516 67790 5568
rect 1012 5466 74980 5488
rect 1012 5414 4210 5466
rect 4262 5414 4274 5466
rect 4326 5414 4338 5466
rect 4390 5414 4402 5466
rect 4454 5414 4466 5466
rect 4518 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 24466 5466
rect 24518 5414 34210 5466
rect 34262 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 44210 5466
rect 44262 5414 44274 5466
rect 44326 5414 44338 5466
rect 44390 5414 44402 5466
rect 44454 5414 44466 5466
rect 44518 5414 54210 5466
rect 54262 5414 54274 5466
rect 54326 5414 54338 5466
rect 54390 5414 54402 5466
rect 54454 5414 54466 5466
rect 54518 5414 64210 5466
rect 64262 5414 64274 5466
rect 64326 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 74210 5466
rect 74262 5414 74274 5466
rect 74326 5414 74338 5466
rect 74390 5414 74402 5466
rect 74454 5414 74466 5466
rect 74518 5414 74980 5466
rect 1012 5392 74980 5414
rect 30116 5324 30880 5352
rect 30116 5293 30144 5324
rect 30101 5287 30159 5293
rect 30101 5253 30113 5287
rect 30147 5253 30159 5287
rect 30101 5247 30159 5253
rect 30742 5244 30748 5296
rect 30800 5244 30806 5296
rect 30852 5284 30880 5324
rect 31018 5312 31024 5364
rect 31076 5312 31082 5364
rect 31386 5312 31392 5364
rect 31444 5352 31450 5364
rect 36446 5352 36452 5364
rect 31444 5324 36452 5352
rect 31444 5312 31450 5324
rect 36446 5312 36452 5324
rect 36504 5312 36510 5364
rect 45278 5352 45284 5364
rect 36556 5324 45284 5352
rect 31110 5284 31116 5296
rect 30852 5256 31116 5284
rect 31110 5244 31116 5256
rect 31168 5244 31174 5296
rect 31202 5244 31208 5296
rect 31260 5284 31266 5296
rect 32398 5284 32404 5296
rect 31260 5256 32404 5284
rect 31260 5244 31266 5256
rect 32398 5244 32404 5256
rect 32456 5244 32462 5296
rect 32582 5244 32588 5296
rect 32640 5284 32646 5296
rect 36556 5284 36584 5324
rect 45278 5312 45284 5324
rect 45336 5312 45342 5364
rect 45370 5312 45376 5364
rect 45428 5352 45434 5364
rect 48498 5352 48504 5364
rect 45428 5324 48504 5352
rect 45428 5312 45434 5324
rect 48498 5312 48504 5324
rect 48556 5312 48562 5364
rect 49053 5355 49111 5361
rect 49053 5321 49065 5355
rect 49099 5352 49111 5355
rect 59078 5352 59084 5364
rect 49099 5324 59084 5352
rect 49099 5321 49111 5324
rect 49053 5315 49111 5321
rect 59078 5312 59084 5324
rect 59136 5312 59142 5364
rect 65978 5312 65984 5364
rect 66036 5352 66042 5364
rect 66254 5352 66260 5364
rect 66036 5324 66260 5352
rect 66036 5312 66042 5324
rect 66254 5312 66260 5324
rect 66312 5312 66318 5364
rect 66530 5312 66536 5364
rect 66588 5312 66594 5364
rect 69198 5312 69204 5364
rect 69256 5312 69262 5364
rect 47210 5284 47216 5296
rect 32640 5256 36584 5284
rect 37384 5256 47216 5284
rect 32640 5244 32646 5256
rect 30377 5219 30435 5225
rect 30377 5185 30389 5219
rect 30423 5216 30435 5219
rect 30558 5216 30564 5228
rect 30423 5188 30564 5216
rect 30423 5185 30435 5188
rect 30377 5179 30435 5185
rect 30558 5176 30564 5188
rect 30616 5216 30622 5228
rect 30926 5216 30932 5228
rect 30616 5188 30932 5216
rect 30616 5176 30622 5188
rect 30926 5176 30932 5188
rect 30984 5176 30990 5228
rect 31294 5176 31300 5228
rect 31352 5216 31358 5228
rect 31481 5219 31539 5225
rect 31481 5216 31493 5219
rect 31352 5188 31493 5216
rect 31352 5176 31358 5188
rect 31481 5185 31493 5188
rect 31527 5216 31539 5219
rect 31662 5216 31668 5228
rect 31527 5188 31668 5216
rect 31527 5185 31539 5188
rect 31481 5179 31539 5185
rect 31662 5176 31668 5188
rect 31720 5176 31726 5228
rect 32490 5176 32496 5228
rect 32548 5176 32554 5228
rect 34606 5176 34612 5228
rect 34664 5216 34670 5228
rect 37384 5216 37412 5256
rect 47210 5244 47216 5256
rect 47268 5244 47274 5296
rect 47302 5244 47308 5296
rect 47360 5244 47366 5296
rect 48133 5287 48191 5293
rect 48133 5253 48145 5287
rect 48179 5284 48191 5287
rect 61746 5284 61752 5296
rect 48179 5256 61752 5284
rect 48179 5253 48191 5256
rect 48133 5247 48191 5253
rect 61746 5244 61752 5256
rect 61804 5244 61810 5296
rect 62117 5287 62175 5293
rect 62117 5253 62129 5287
rect 62163 5284 62175 5287
rect 62298 5284 62304 5296
rect 62163 5256 62304 5284
rect 62163 5253 62175 5256
rect 62117 5247 62175 5253
rect 62298 5244 62304 5256
rect 62356 5244 62362 5296
rect 62390 5244 62396 5296
rect 62448 5284 62454 5296
rect 63862 5284 63868 5296
rect 62448 5256 63868 5284
rect 62448 5244 62454 5256
rect 63862 5244 63868 5256
rect 63920 5244 63926 5296
rect 65334 5216 65340 5228
rect 34664 5188 37412 5216
rect 41386 5188 45692 5216
rect 34664 5176 34670 5188
rect 32306 5108 32312 5160
rect 32364 5108 32370 5160
rect 32398 5108 32404 5160
rect 32456 5148 32462 5160
rect 41386 5148 41414 5188
rect 32456 5120 41414 5148
rect 32456 5108 32462 5120
rect 43898 5108 43904 5160
rect 43956 5148 43962 5160
rect 44637 5151 44695 5157
rect 44637 5148 44649 5151
rect 43956 5120 44649 5148
rect 43956 5108 43962 5120
rect 44637 5117 44649 5120
rect 44683 5148 44695 5151
rect 44821 5151 44879 5157
rect 44821 5148 44833 5151
rect 44683 5120 44833 5148
rect 44683 5117 44695 5120
rect 44637 5111 44695 5117
rect 44821 5117 44833 5120
rect 44867 5117 44879 5151
rect 44821 5111 44879 5117
rect 44910 5108 44916 5160
rect 44968 5148 44974 5160
rect 45554 5148 45560 5160
rect 44968 5120 45560 5148
rect 44968 5108 44974 5120
rect 45554 5108 45560 5120
rect 45612 5108 45618 5160
rect 45664 5148 45692 5188
rect 47504 5188 65340 5216
rect 47504 5148 47532 5188
rect 65334 5176 65340 5188
rect 65392 5176 65398 5228
rect 45664 5120 47532 5148
rect 47578 5108 47584 5160
rect 47636 5148 47642 5160
rect 48225 5151 48283 5157
rect 48225 5148 48237 5151
rect 47636 5120 48237 5148
rect 47636 5108 47642 5120
rect 48225 5117 48237 5120
rect 48271 5117 48283 5151
rect 48225 5111 48283 5117
rect 48406 5108 48412 5160
rect 48464 5108 48470 5160
rect 48498 5108 48504 5160
rect 48556 5148 48562 5160
rect 50525 5151 50583 5157
rect 50525 5148 50537 5151
rect 48556 5120 50537 5148
rect 48556 5108 48562 5120
rect 50525 5117 50537 5120
rect 50571 5117 50583 5151
rect 50525 5111 50583 5117
rect 52454 5108 52460 5160
rect 52512 5148 52518 5160
rect 54297 5151 54355 5157
rect 54297 5148 54309 5151
rect 52512 5120 54309 5148
rect 52512 5108 52518 5120
rect 54297 5117 54309 5120
rect 54343 5117 54355 5151
rect 60274 5148 60280 5160
rect 54297 5111 54355 5117
rect 54404 5120 60280 5148
rect 29914 5040 29920 5092
rect 29972 5040 29978 5092
rect 32214 5040 32220 5092
rect 32272 5080 32278 5092
rect 32272 5052 44036 5080
rect 32272 5040 32278 5052
rect 30834 4972 30840 5024
rect 30892 5012 30898 5024
rect 31386 5012 31392 5024
rect 30892 4984 31392 5012
rect 30892 4972 30898 4984
rect 31386 4972 31392 4984
rect 31444 4972 31450 5024
rect 34698 4972 34704 5024
rect 34756 4972 34762 5024
rect 35158 4972 35164 5024
rect 35216 5012 35222 5024
rect 35526 5012 35532 5024
rect 35216 4984 35532 5012
rect 35216 4972 35222 4984
rect 35526 4972 35532 4984
rect 35584 4972 35590 5024
rect 36446 4972 36452 5024
rect 36504 5012 36510 5024
rect 43898 5012 43904 5024
rect 36504 4984 43904 5012
rect 36504 4972 36510 4984
rect 43898 4972 43904 4984
rect 43956 4972 43962 5024
rect 44008 5012 44036 5052
rect 45462 5040 45468 5092
rect 45520 5040 45526 5092
rect 54404 5080 54432 5120
rect 60274 5108 60280 5120
rect 60332 5108 60338 5160
rect 62758 5148 62764 5160
rect 61028 5120 62764 5148
rect 61028 5080 61056 5120
rect 62758 5108 62764 5120
rect 62816 5108 62822 5160
rect 45572 5052 54432 5080
rect 54864 5052 61056 5080
rect 45572 5012 45600 5052
rect 44008 4984 45600 5012
rect 45738 4972 45744 5024
rect 45796 5012 45802 5024
rect 49050 5012 49056 5024
rect 45796 4984 49056 5012
rect 45796 4972 45802 4984
rect 49050 4972 49056 4984
rect 49108 4972 49114 5024
rect 51169 5015 51227 5021
rect 51169 4981 51181 5015
rect 51215 5012 51227 5015
rect 54864 5012 54892 5052
rect 61102 5040 61108 5092
rect 61160 5080 61166 5092
rect 63770 5080 63776 5092
rect 61160 5052 63776 5080
rect 61160 5040 61166 5052
rect 63770 5040 63776 5052
rect 63828 5040 63834 5092
rect 51215 4984 54892 5012
rect 54941 5015 54999 5021
rect 51215 4981 51227 4984
rect 51169 4975 51227 4981
rect 54941 4981 54953 5015
rect 54987 5012 54999 5015
rect 58894 5012 58900 5024
rect 54987 4984 58900 5012
rect 54987 4981 54999 4984
rect 54941 4975 54999 4981
rect 58894 4972 58900 4984
rect 58952 4972 58958 5024
rect 59170 4972 59176 5024
rect 59228 4972 59234 5024
rect 60553 5015 60611 5021
rect 60553 4981 60565 5015
rect 60599 5012 60611 5015
rect 60734 5012 60740 5024
rect 60599 4984 60740 5012
rect 60599 4981 60611 4984
rect 60553 4975 60611 4981
rect 60734 4972 60740 4984
rect 60792 4972 60798 5024
rect 63586 4972 63592 5024
rect 63644 4972 63650 5024
rect 1012 4922 74980 4944
rect 1012 4870 1858 4922
rect 1910 4870 1922 4922
rect 1974 4870 1986 4922
rect 2038 4870 2050 4922
rect 2102 4870 2114 4922
rect 2166 4870 11858 4922
rect 11910 4870 11922 4922
rect 11974 4870 11986 4922
rect 12038 4870 12050 4922
rect 12102 4870 12114 4922
rect 12166 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 21986 4922
rect 22038 4870 22050 4922
rect 22102 4870 22114 4922
rect 22166 4870 31858 4922
rect 31910 4870 31922 4922
rect 31974 4870 31986 4922
rect 32038 4870 32050 4922
rect 32102 4870 32114 4922
rect 32166 4870 41858 4922
rect 41910 4870 41922 4922
rect 41974 4870 41986 4922
rect 42038 4870 42050 4922
rect 42102 4870 42114 4922
rect 42166 4870 51858 4922
rect 51910 4870 51922 4922
rect 51974 4870 51986 4922
rect 52038 4870 52050 4922
rect 52102 4870 52114 4922
rect 52166 4870 61858 4922
rect 61910 4870 61922 4922
rect 61974 4870 61986 4922
rect 62038 4870 62050 4922
rect 62102 4870 62114 4922
rect 62166 4870 71858 4922
rect 71910 4870 71922 4922
rect 71974 4870 71986 4922
rect 72038 4870 72050 4922
rect 72102 4870 72114 4922
rect 72166 4870 74980 4922
rect 1012 4848 74980 4870
rect 30193 4811 30251 4817
rect 30193 4777 30205 4811
rect 30239 4808 30251 4811
rect 31202 4808 31208 4820
rect 30239 4780 31208 4808
rect 30239 4777 30251 4780
rect 30193 4771 30251 4777
rect 31202 4768 31208 4780
rect 31260 4768 31266 4820
rect 31573 4811 31631 4817
rect 31573 4777 31585 4811
rect 31619 4808 31631 4811
rect 32398 4808 32404 4820
rect 31619 4780 32404 4808
rect 31619 4777 31631 4780
rect 31573 4771 31631 4777
rect 32398 4768 32404 4780
rect 32456 4768 32462 4820
rect 34054 4808 34060 4820
rect 32508 4780 34060 4808
rect 32306 4740 32312 4752
rect 29104 4712 32312 4740
rect 29104 4613 29132 4712
rect 32306 4700 32312 4712
rect 32364 4700 32370 4752
rect 29825 4675 29883 4681
rect 29825 4641 29837 4675
rect 29871 4672 29883 4675
rect 29914 4672 29920 4684
rect 29871 4644 29920 4672
rect 29871 4641 29883 4644
rect 29825 4635 29883 4641
rect 29914 4632 29920 4644
rect 29972 4632 29978 4684
rect 30009 4675 30067 4681
rect 30009 4641 30021 4675
rect 30055 4672 30067 4675
rect 32508 4672 32536 4780
rect 34054 4768 34060 4780
rect 34112 4768 34118 4820
rect 35713 4811 35771 4817
rect 34532 4780 34744 4808
rect 34532 4740 34560 4780
rect 32600 4712 34560 4740
rect 34609 4743 34667 4749
rect 32600 4681 32628 4712
rect 34609 4709 34621 4743
rect 34655 4709 34667 4743
rect 34716 4740 34744 4780
rect 35713 4777 35725 4811
rect 35759 4808 35771 4811
rect 35759 4780 45416 4808
rect 35759 4777 35771 4780
rect 35713 4771 35771 4777
rect 45388 4740 45416 4780
rect 45462 4768 45468 4820
rect 45520 4808 45526 4820
rect 60458 4808 60464 4820
rect 45520 4780 60464 4808
rect 45520 4768 45526 4780
rect 60458 4768 60464 4780
rect 60516 4768 60522 4820
rect 62117 4811 62175 4817
rect 62117 4777 62129 4811
rect 62163 4808 62175 4811
rect 62298 4808 62304 4820
rect 62163 4780 62304 4808
rect 62163 4777 62175 4780
rect 62117 4771 62175 4777
rect 62298 4768 62304 4780
rect 62356 4768 62362 4820
rect 66530 4768 66536 4820
rect 66588 4768 66594 4820
rect 69198 4768 69204 4820
rect 69256 4768 69262 4820
rect 45738 4740 45744 4752
rect 34716 4712 41414 4740
rect 45388 4712 45744 4740
rect 34609 4703 34667 4709
rect 30055 4644 32536 4672
rect 32585 4675 32643 4681
rect 30055 4641 30067 4644
rect 30009 4635 30067 4641
rect 32585 4641 32597 4675
rect 32631 4641 32643 4675
rect 32585 4635 32643 4641
rect 33962 4632 33968 4684
rect 34020 4672 34026 4684
rect 34624 4672 34652 4703
rect 34020 4644 34652 4672
rect 34768 4675 34826 4681
rect 34020 4632 34026 4644
rect 34768 4641 34780 4675
rect 34814 4672 34826 4675
rect 34974 4672 34980 4684
rect 34814 4644 34980 4672
rect 34814 4641 34826 4644
rect 34768 4635 34826 4641
rect 34974 4632 34980 4644
rect 35032 4632 35038 4684
rect 35253 4675 35311 4681
rect 35253 4641 35265 4675
rect 35299 4672 35311 4675
rect 35299 4644 35480 4672
rect 35299 4641 35311 4644
rect 35253 4635 35311 4641
rect 28905 4607 28963 4613
rect 28905 4573 28917 4607
rect 28951 4573 28963 4607
rect 28905 4567 28963 4573
rect 29089 4607 29147 4613
rect 29089 4573 29101 4607
rect 29135 4573 29147 4607
rect 29089 4567 29147 4573
rect 29273 4607 29331 4613
rect 29273 4573 29285 4607
rect 29319 4604 29331 4607
rect 29362 4604 29368 4616
rect 29319 4576 29368 4604
rect 29319 4573 29331 4576
rect 29273 4567 29331 4573
rect 28629 4539 28687 4545
rect 28629 4505 28641 4539
rect 28675 4505 28687 4539
rect 28920 4536 28948 4567
rect 29362 4564 29368 4576
rect 29420 4604 29426 4616
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 29420 4576 29561 4604
rect 29420 4564 29426 4576
rect 29549 4573 29561 4576
rect 29595 4604 29607 4607
rect 30926 4604 30932 4616
rect 29595 4576 30932 4604
rect 29595 4573 29607 4576
rect 29549 4567 29607 4573
rect 30926 4564 30932 4576
rect 30984 4564 30990 4616
rect 32766 4564 32772 4616
rect 32824 4564 32830 4616
rect 32858 4564 32864 4616
rect 32916 4604 32922 4616
rect 34241 4607 34299 4613
rect 32916 4576 34008 4604
rect 32916 4564 32922 4576
rect 33980 4548 34008 4576
rect 34241 4573 34253 4607
rect 34287 4604 34299 4607
rect 34606 4604 34612 4616
rect 34287 4576 34612 4604
rect 34287 4573 34299 4576
rect 34241 4567 34299 4573
rect 34606 4564 34612 4576
rect 34664 4564 34670 4616
rect 34885 4607 34943 4613
rect 34885 4604 34897 4607
rect 34808 4576 34897 4604
rect 29454 4536 29460 4548
rect 28920 4508 29460 4536
rect 28629 4499 28687 4505
rect 28644 4468 28672 4499
rect 29454 4496 29460 4508
rect 29512 4496 29518 4548
rect 30466 4496 30472 4548
rect 30524 4496 30530 4548
rect 30742 4496 30748 4548
rect 30800 4496 30806 4548
rect 31110 4496 31116 4548
rect 31168 4536 31174 4548
rect 31414 4539 31472 4545
rect 31414 4536 31426 4539
rect 31168 4508 31426 4536
rect 31168 4496 31174 4508
rect 31414 4505 31426 4508
rect 31460 4505 31472 4539
rect 31414 4499 31472 4505
rect 33870 4496 33876 4548
rect 33928 4496 33934 4548
rect 33962 4496 33968 4548
rect 34020 4496 34026 4548
rect 34808 4536 34836 4576
rect 34885 4573 34897 4576
rect 34931 4604 34943 4607
rect 35158 4604 35164 4616
rect 34931 4576 35164 4604
rect 34931 4573 34943 4576
rect 34885 4567 34943 4573
rect 35158 4564 35164 4576
rect 35216 4564 35222 4616
rect 35452 4604 35480 4644
rect 36262 4632 36268 4684
rect 36320 4672 36326 4684
rect 40034 4672 40040 4684
rect 36320 4644 40040 4672
rect 36320 4632 36326 4644
rect 40034 4632 40040 4644
rect 40092 4632 40098 4684
rect 41386 4672 41414 4712
rect 45738 4700 45744 4712
rect 45796 4700 45802 4752
rect 59262 4740 59268 4752
rect 46768 4712 59268 4740
rect 46566 4672 46572 4684
rect 41386 4644 46572 4672
rect 46566 4632 46572 4644
rect 46624 4632 46630 4684
rect 46768 4681 46796 4712
rect 59262 4700 59268 4712
rect 59320 4700 59326 4752
rect 61194 4700 61200 4752
rect 61252 4700 61258 4752
rect 63586 4700 63592 4752
rect 63644 4740 63650 4752
rect 63954 4740 63960 4752
rect 63644 4712 63960 4740
rect 63644 4700 63650 4712
rect 63954 4700 63960 4712
rect 64012 4700 64018 4752
rect 46753 4675 46811 4681
rect 46753 4641 46765 4675
rect 46799 4641 46811 4675
rect 46753 4635 46811 4641
rect 46934 4632 46940 4684
rect 46992 4672 46998 4684
rect 59354 4672 59360 4684
rect 46992 4644 59360 4672
rect 46992 4632 46998 4644
rect 59354 4632 59360 4644
rect 59412 4632 59418 4684
rect 35710 4604 35716 4616
rect 35452 4576 35716 4604
rect 35710 4564 35716 4576
rect 35768 4564 35774 4616
rect 36170 4564 36176 4616
rect 36228 4604 36234 4616
rect 36228 4576 41414 4604
rect 36228 4564 36234 4576
rect 34072 4508 34836 4536
rect 29822 4468 29828 4480
rect 28644 4440 29828 4468
rect 29822 4428 29828 4440
rect 29880 4428 29886 4480
rect 29917 4471 29975 4477
rect 29917 4437 29929 4471
rect 29963 4468 29975 4471
rect 30650 4468 30656 4480
rect 29963 4440 30656 4468
rect 29963 4437 29975 4440
rect 29917 4431 29975 4437
rect 30650 4428 30656 4440
rect 30708 4428 30714 4480
rect 31018 4428 31024 4480
rect 31076 4468 31082 4480
rect 31205 4471 31263 4477
rect 31205 4468 31217 4471
rect 31076 4440 31217 4468
rect 31076 4428 31082 4440
rect 31205 4437 31217 4440
rect 31251 4437 31263 4471
rect 31205 4431 31263 4437
rect 31294 4428 31300 4480
rect 31352 4428 31358 4480
rect 32125 4471 32183 4477
rect 32125 4437 32137 4471
rect 32171 4468 32183 4471
rect 32950 4468 32956 4480
rect 32171 4440 32956 4468
rect 32171 4437 32183 4440
rect 32125 4431 32183 4437
rect 32950 4428 32956 4440
rect 33008 4428 33014 4480
rect 33594 4428 33600 4480
rect 33652 4468 33658 4480
rect 34072 4468 34100 4508
rect 35066 4496 35072 4548
rect 35124 4536 35130 4548
rect 35437 4539 35495 4545
rect 35437 4536 35449 4539
rect 35124 4508 35449 4536
rect 35124 4496 35130 4508
rect 35437 4505 35449 4508
rect 35483 4505 35495 4539
rect 41386 4536 41414 4576
rect 44726 4564 44732 4616
rect 44784 4604 44790 4616
rect 45557 4607 45615 4613
rect 45557 4604 45569 4607
rect 44784 4576 45569 4604
rect 44784 4564 44790 4576
rect 45557 4573 45569 4576
rect 45603 4573 45615 4607
rect 45557 4567 45615 4573
rect 45664 4576 46612 4604
rect 45664 4536 45692 4576
rect 41386 4508 45692 4536
rect 46584 4536 46612 4576
rect 46842 4564 46848 4616
rect 46900 4604 46906 4616
rect 47489 4607 47547 4613
rect 47489 4604 47501 4607
rect 46900 4576 47501 4604
rect 46900 4564 46906 4576
rect 47489 4573 47501 4576
rect 47535 4573 47547 4607
rect 59998 4604 60004 4616
rect 47489 4567 47547 4573
rect 47596 4576 60004 4604
rect 47596 4536 47624 4576
rect 59998 4564 60004 4576
rect 60056 4564 60062 4616
rect 60553 4607 60611 4613
rect 60553 4573 60565 4607
rect 60599 4604 60611 4607
rect 60642 4604 60648 4616
rect 60599 4576 60648 4604
rect 60599 4573 60611 4576
rect 60553 4567 60611 4573
rect 60642 4564 60648 4576
rect 60700 4564 60706 4616
rect 46584 4508 47624 4536
rect 48685 4539 48743 4545
rect 35437 4499 35495 4505
rect 48685 4505 48697 4539
rect 48731 4536 48743 4539
rect 53742 4536 53748 4548
rect 48731 4508 53748 4536
rect 48731 4505 48743 4508
rect 48685 4499 48743 4505
rect 53742 4496 53748 4508
rect 53800 4496 53806 4548
rect 59538 4536 59544 4548
rect 53944 4508 59544 4536
rect 33652 4440 34100 4468
rect 34977 4471 35035 4477
rect 33652 4428 33658 4440
rect 34977 4437 34989 4471
rect 35023 4468 35035 4471
rect 35158 4468 35164 4480
rect 35023 4440 35164 4468
rect 35023 4437 35035 4440
rect 34977 4431 35035 4437
rect 35158 4428 35164 4440
rect 35216 4428 35222 4480
rect 35618 4428 35624 4480
rect 35676 4468 35682 4480
rect 53944 4468 53972 4508
rect 59538 4496 59544 4508
rect 59596 4496 59602 4548
rect 60734 4496 60740 4548
rect 60792 4536 60798 4548
rect 61038 4539 61096 4545
rect 61038 4536 61050 4539
rect 60792 4508 61050 4536
rect 60792 4496 60798 4508
rect 61038 4505 61050 4508
rect 61084 4505 61096 4539
rect 61038 4499 61096 4505
rect 61470 4496 61476 4548
rect 61528 4536 61534 4548
rect 65058 4536 65064 4548
rect 61528 4508 65064 4536
rect 61528 4496 61534 4508
rect 65058 4496 65064 4508
rect 65116 4496 65122 4548
rect 35676 4440 53972 4468
rect 35676 4428 35682 4440
rect 59170 4428 59176 4480
rect 59228 4428 59234 4480
rect 59354 4428 59360 4480
rect 59412 4468 59418 4480
rect 60826 4468 60832 4480
rect 59412 4440 60832 4468
rect 59412 4428 59418 4440
rect 60826 4428 60832 4440
rect 60884 4428 60890 4480
rect 60918 4428 60924 4480
rect 60976 4428 60982 4480
rect 62758 4428 62764 4480
rect 62816 4468 62822 4480
rect 70118 4468 70124 4480
rect 62816 4440 70124 4468
rect 62816 4428 62822 4440
rect 70118 4428 70124 4440
rect 70176 4428 70182 4480
rect 1012 4378 74980 4400
rect 1012 4326 4210 4378
rect 4262 4326 4274 4378
rect 4326 4326 4338 4378
rect 4390 4326 4402 4378
rect 4454 4326 4466 4378
rect 4518 4326 14210 4378
rect 14262 4326 14274 4378
rect 14326 4326 14338 4378
rect 14390 4326 14402 4378
rect 14454 4326 14466 4378
rect 14518 4326 24210 4378
rect 24262 4326 24274 4378
rect 24326 4326 24338 4378
rect 24390 4326 24402 4378
rect 24454 4326 24466 4378
rect 24518 4326 34210 4378
rect 34262 4326 34274 4378
rect 34326 4326 34338 4378
rect 34390 4326 34402 4378
rect 34454 4326 34466 4378
rect 34518 4326 44210 4378
rect 44262 4326 44274 4378
rect 44326 4326 44338 4378
rect 44390 4326 44402 4378
rect 44454 4326 44466 4378
rect 44518 4326 54210 4378
rect 54262 4326 54274 4378
rect 54326 4326 54338 4378
rect 54390 4326 54402 4378
rect 54454 4326 54466 4378
rect 54518 4326 64210 4378
rect 64262 4326 64274 4378
rect 64326 4326 64338 4378
rect 64390 4326 64402 4378
rect 64454 4326 64466 4378
rect 64518 4326 74210 4378
rect 74262 4326 74274 4378
rect 74326 4326 74338 4378
rect 74390 4326 74402 4378
rect 74454 4326 74466 4378
rect 74518 4326 74980 4378
rect 1012 4304 74980 4326
rect 29733 4267 29791 4273
rect 29733 4233 29745 4267
rect 29779 4264 29791 4267
rect 30650 4264 30656 4276
rect 29779 4236 30656 4264
rect 29779 4233 29791 4236
rect 29733 4227 29791 4233
rect 30650 4224 30656 4236
rect 30708 4264 30714 4276
rect 30745 4267 30803 4273
rect 30745 4264 30757 4267
rect 30708 4236 30757 4264
rect 30708 4224 30714 4236
rect 30745 4233 30757 4236
rect 30791 4264 30803 4267
rect 31294 4264 31300 4276
rect 30791 4236 31300 4264
rect 30791 4233 30803 4236
rect 30745 4227 30803 4233
rect 31294 4224 31300 4236
rect 31352 4264 31358 4276
rect 31573 4267 31631 4273
rect 31573 4264 31585 4267
rect 31352 4236 31585 4264
rect 31352 4224 31358 4236
rect 31573 4233 31585 4236
rect 31619 4264 31631 4267
rect 32493 4267 32551 4273
rect 32493 4264 32505 4267
rect 31619 4236 32505 4264
rect 31619 4233 31631 4236
rect 31573 4227 31631 4233
rect 32493 4233 32505 4236
rect 32539 4264 32551 4267
rect 33594 4264 33600 4276
rect 32539 4236 33600 4264
rect 32539 4233 32551 4236
rect 32493 4227 32551 4233
rect 33594 4224 33600 4236
rect 33652 4264 33658 4276
rect 33689 4267 33747 4273
rect 33689 4264 33701 4267
rect 33652 4236 33701 4264
rect 33652 4224 33658 4236
rect 33689 4233 33701 4236
rect 33735 4233 33747 4267
rect 33689 4227 33747 4233
rect 33781 4267 33839 4273
rect 33781 4233 33793 4267
rect 33827 4264 33839 4267
rect 34054 4264 34060 4276
rect 33827 4236 34060 4264
rect 33827 4233 33839 4236
rect 33781 4227 33839 4233
rect 34054 4224 34060 4236
rect 34112 4224 34118 4276
rect 34333 4267 34391 4273
rect 34333 4264 34345 4267
rect 34164 4236 34345 4264
rect 29362 4156 29368 4208
rect 29420 4156 29426 4208
rect 29641 4199 29699 4205
rect 29641 4165 29653 4199
rect 29687 4196 29699 4199
rect 29914 4196 29920 4208
rect 29687 4168 29920 4196
rect 29687 4165 29699 4168
rect 29641 4159 29699 4165
rect 29914 4156 29920 4168
rect 29972 4156 29978 4208
rect 30466 4156 30472 4208
rect 30524 4196 30530 4208
rect 30837 4199 30895 4205
rect 30837 4196 30849 4199
rect 30524 4168 30849 4196
rect 30524 4156 30530 4168
rect 30837 4165 30849 4168
rect 30883 4165 30895 4199
rect 30837 4159 30895 4165
rect 32610 4199 32668 4205
rect 32610 4165 32622 4199
rect 32656 4196 32668 4199
rect 32950 4196 32956 4208
rect 32656 4168 32956 4196
rect 32656 4165 32668 4168
rect 32610 4159 32668 4165
rect 32950 4156 32956 4168
rect 33008 4156 33014 4208
rect 33962 4156 33968 4208
rect 34020 4196 34026 4208
rect 34164 4196 34192 4236
rect 34333 4233 34345 4236
rect 34379 4233 34391 4267
rect 34333 4227 34391 4233
rect 34609 4267 34667 4273
rect 34609 4233 34621 4267
rect 34655 4264 34667 4267
rect 34882 4264 34888 4276
rect 34655 4236 34888 4264
rect 34655 4233 34667 4236
rect 34609 4227 34667 4233
rect 34882 4224 34888 4236
rect 34940 4224 34946 4276
rect 34974 4224 34980 4276
rect 35032 4264 35038 4276
rect 35069 4267 35127 4273
rect 35069 4264 35081 4267
rect 35032 4236 35081 4264
rect 35032 4224 35038 4236
rect 35069 4233 35081 4236
rect 35115 4233 35127 4267
rect 35069 4227 35127 4233
rect 35342 4224 35348 4276
rect 35400 4224 35406 4276
rect 35802 4224 35808 4276
rect 35860 4264 35866 4276
rect 35860 4236 40724 4264
rect 35860 4224 35866 4236
rect 34020 4168 34192 4196
rect 34020 4156 34026 4168
rect 34698 4156 34704 4208
rect 34756 4156 34762 4208
rect 35228 4199 35286 4205
rect 35228 4165 35240 4199
rect 35274 4165 35286 4199
rect 35228 4159 35286 4165
rect 30285 4131 30343 4137
rect 30285 4097 30297 4131
rect 30331 4128 30343 4131
rect 30484 4128 30512 4156
rect 30926 4128 30932 4140
rect 30331 4100 30512 4128
rect 30576 4100 30932 4128
rect 30331 4097 30343 4100
rect 30285 4091 30343 4097
rect 28074 4020 28080 4072
rect 28132 4020 28138 4072
rect 28994 4020 29000 4072
rect 29052 4060 29058 4072
rect 29181 4063 29239 4069
rect 29181 4060 29193 4063
rect 29052 4032 29193 4060
rect 29052 4020 29058 4032
rect 29181 4029 29193 4032
rect 29227 4029 29239 4063
rect 29181 4023 29239 4029
rect 29822 4020 29828 4072
rect 29880 4020 29886 4072
rect 30377 4063 30435 4069
rect 30377 4029 30389 4063
rect 30423 4060 30435 4063
rect 30576 4060 30604 4100
rect 30926 4088 30932 4100
rect 30984 4128 30990 4140
rect 31205 4131 31263 4137
rect 31205 4128 31217 4131
rect 30984 4100 31217 4128
rect 30984 4088 30990 4100
rect 31205 4097 31217 4100
rect 31251 4128 31263 4131
rect 32125 4131 32183 4137
rect 32125 4128 32137 4131
rect 31251 4100 32137 4128
rect 31251 4097 31263 4100
rect 31205 4091 31263 4097
rect 32125 4097 32137 4100
rect 32171 4128 32183 4131
rect 35243 4128 35271 4159
rect 35434 4156 35440 4208
rect 35492 4156 35498 4208
rect 35894 4156 35900 4208
rect 35952 4196 35958 4208
rect 40696 4196 40724 4236
rect 40770 4224 40776 4276
rect 40828 4264 40834 4276
rect 46937 4267 46995 4273
rect 46937 4264 46949 4267
rect 40828 4236 46949 4264
rect 40828 4224 40834 4236
rect 46937 4233 46949 4236
rect 46983 4264 46995 4267
rect 48501 4267 48559 4273
rect 48501 4264 48513 4267
rect 46983 4236 48513 4264
rect 46983 4233 46995 4236
rect 46937 4227 46995 4233
rect 48501 4233 48513 4236
rect 48547 4264 48559 4267
rect 50157 4267 50215 4273
rect 50157 4264 50169 4267
rect 48547 4236 50169 4264
rect 48547 4233 48559 4236
rect 48501 4227 48559 4233
rect 50157 4233 50169 4236
rect 50203 4264 50215 4267
rect 51721 4267 51779 4273
rect 51721 4264 51733 4267
rect 50203 4236 51733 4264
rect 50203 4233 50215 4236
rect 50157 4227 50215 4233
rect 51721 4233 51733 4236
rect 51767 4264 51779 4267
rect 53193 4267 53251 4273
rect 53193 4264 53205 4267
rect 51767 4236 53205 4264
rect 51767 4233 51779 4236
rect 51721 4227 51779 4233
rect 53193 4233 53205 4236
rect 53239 4264 53251 4267
rect 54849 4267 54907 4273
rect 54849 4264 54861 4267
rect 53239 4236 54861 4264
rect 53239 4233 53251 4236
rect 53193 4227 53251 4233
rect 54849 4233 54861 4236
rect 54895 4264 54907 4267
rect 56321 4267 56379 4273
rect 56321 4264 56333 4267
rect 54895 4236 56333 4264
rect 54895 4233 54907 4236
rect 54849 4227 54907 4233
rect 56321 4233 56333 4236
rect 56367 4264 56379 4267
rect 58069 4267 58127 4273
rect 58069 4264 58081 4267
rect 56367 4236 58081 4264
rect 56367 4233 56379 4236
rect 56321 4227 56379 4233
rect 58069 4233 58081 4236
rect 58115 4264 58127 4267
rect 59354 4264 59360 4276
rect 58115 4236 59360 4264
rect 58115 4233 58127 4236
rect 58069 4227 58127 4233
rect 59354 4224 59360 4236
rect 59412 4224 59418 4276
rect 60550 4224 60556 4276
rect 60608 4264 60614 4276
rect 60645 4267 60703 4273
rect 60645 4264 60657 4267
rect 60608 4236 60657 4264
rect 60608 4224 60614 4236
rect 60645 4233 60657 4236
rect 60691 4264 60703 4267
rect 60734 4264 60740 4276
rect 60691 4236 60740 4264
rect 60691 4233 60703 4236
rect 60645 4227 60703 4233
rect 60734 4224 60740 4236
rect 60792 4224 60798 4276
rect 60826 4224 60832 4276
rect 60884 4264 60890 4276
rect 62301 4267 62359 4273
rect 62301 4264 62313 4267
rect 60884 4236 62313 4264
rect 60884 4224 60890 4236
rect 62301 4233 62313 4236
rect 62347 4264 62359 4267
rect 63773 4267 63831 4273
rect 63773 4264 63785 4267
rect 62347 4236 63785 4264
rect 62347 4233 62359 4236
rect 62301 4227 62359 4233
rect 63773 4233 63785 4236
rect 63819 4233 63831 4267
rect 63773 4227 63831 4233
rect 65242 4224 65248 4276
rect 65300 4264 65306 4276
rect 66717 4267 66775 4273
rect 66717 4264 66729 4267
rect 65300 4236 66729 4264
rect 65300 4224 65306 4236
rect 66717 4233 66729 4236
rect 66763 4264 66775 4267
rect 68373 4267 68431 4273
rect 68373 4264 68385 4267
rect 66763 4236 68385 4264
rect 66763 4233 66775 4236
rect 66717 4227 66775 4233
rect 68373 4233 68385 4236
rect 68419 4264 68431 4267
rect 69477 4267 69535 4273
rect 69477 4264 69489 4267
rect 68419 4236 69489 4264
rect 68419 4233 68431 4236
rect 68373 4227 68431 4233
rect 69477 4233 69489 4236
rect 69523 4233 69535 4267
rect 69477 4227 69535 4233
rect 47029 4199 47087 4205
rect 47029 4196 47041 4199
rect 35952 4168 40632 4196
rect 35952 4156 35958 4168
rect 35526 4128 35532 4140
rect 32171 4100 32996 4128
rect 35243 4100 35532 4128
rect 32171 4097 32183 4100
rect 32125 4091 32183 4097
rect 32968 4072 32996 4100
rect 35526 4088 35532 4100
rect 35584 4088 35590 4140
rect 35710 4088 35716 4140
rect 35768 4088 35774 4140
rect 35802 4088 35808 4140
rect 35860 4128 35866 4140
rect 35989 4131 36047 4137
rect 35989 4128 36001 4131
rect 35860 4100 36001 4128
rect 35860 4088 35866 4100
rect 35989 4097 36001 4100
rect 36035 4097 36047 4131
rect 35989 4091 36047 4097
rect 36630 4088 36636 4140
rect 36688 4088 36694 4140
rect 30423 4032 30604 4060
rect 30423 4029 30435 4032
rect 30377 4023 30435 4029
rect 30650 4020 30656 4072
rect 30708 4060 30714 4072
rect 31018 4060 31024 4072
rect 30708 4032 31024 4060
rect 30708 4020 30714 4032
rect 31018 4020 31024 4032
rect 31076 4060 31082 4072
rect 31481 4063 31539 4069
rect 31481 4060 31493 4063
rect 31076 4032 31493 4060
rect 31076 4020 31082 4032
rect 31481 4029 31493 4032
rect 31527 4029 31539 4063
rect 31481 4023 31539 4029
rect 31662 4020 31668 4072
rect 31720 4069 31726 4072
rect 31720 4063 31748 4069
rect 31736 4029 31748 4063
rect 31720 4023 31748 4029
rect 31720 4020 31726 4023
rect 32306 4020 32312 4072
rect 32364 4060 32370 4072
rect 32401 4063 32459 4069
rect 32401 4060 32413 4063
rect 32364 4032 32413 4060
rect 32364 4020 32370 4032
rect 32401 4029 32413 4032
rect 32447 4029 32459 4063
rect 32401 4023 32459 4029
rect 32950 4020 32956 4072
rect 33008 4020 33014 4072
rect 33318 4020 33324 4072
rect 33376 4060 33382 4072
rect 33572 4063 33630 4069
rect 33572 4060 33584 4063
rect 33376 4032 33584 4060
rect 33376 4020 33382 4032
rect 33572 4029 33584 4032
rect 33618 4060 33630 4063
rect 33686 4060 33692 4072
rect 33618 4032 33692 4060
rect 33618 4029 33630 4032
rect 33572 4023 33630 4029
rect 33686 4020 33692 4032
rect 33744 4020 33750 4072
rect 34054 4020 34060 4072
rect 34112 4020 34118 4072
rect 34241 4063 34299 4069
rect 34241 4029 34253 4063
rect 34287 4060 34299 4063
rect 34492 4063 34550 4069
rect 34492 4060 34504 4063
rect 34287 4032 34504 4060
rect 34287 4029 34299 4032
rect 34241 4023 34299 4029
rect 34492 4029 34504 4032
rect 34538 4060 34550 4063
rect 34790 4060 34796 4072
rect 34538 4032 34796 4060
rect 34538 4029 34550 4032
rect 34492 4023 34550 4029
rect 34790 4020 34796 4032
rect 34848 4020 34854 4072
rect 34977 4063 35035 4069
rect 34977 4029 34989 4063
rect 35023 4060 35035 4063
rect 35023 4032 35204 4060
rect 35023 4029 35035 4032
rect 34977 4023 35035 4029
rect 30009 3995 30067 4001
rect 30009 3961 30021 3995
rect 30055 3992 30067 3995
rect 32582 3992 32588 4004
rect 30055 3964 32588 3992
rect 30055 3961 30067 3964
rect 30009 3955 30067 3961
rect 32582 3952 32588 3964
rect 32640 3952 32646 4004
rect 34992 3992 35020 4023
rect 32692 3964 35020 3992
rect 35176 3992 35204 4032
rect 36262 4020 36268 4072
rect 36320 4020 36326 4072
rect 40218 4020 40224 4072
rect 40276 4020 40282 4072
rect 40604 4060 40632 4168
rect 40696 4168 47041 4196
rect 40696 4137 40724 4168
rect 47029 4165 47041 4168
rect 47075 4196 47087 4199
rect 48593 4199 48651 4205
rect 48593 4196 48605 4199
rect 47075 4168 48605 4196
rect 47075 4165 47087 4168
rect 47029 4159 47087 4165
rect 48593 4165 48605 4168
rect 48639 4196 48651 4199
rect 50249 4199 50307 4205
rect 50249 4196 50261 4199
rect 48639 4168 50261 4196
rect 48639 4165 48651 4168
rect 48593 4159 48651 4165
rect 50249 4165 50261 4168
rect 50295 4196 50307 4199
rect 51813 4199 51871 4205
rect 51813 4196 51825 4199
rect 50295 4168 51825 4196
rect 50295 4165 50307 4168
rect 50249 4159 50307 4165
rect 51813 4165 51825 4168
rect 51859 4196 51871 4199
rect 53285 4199 53343 4205
rect 53285 4196 53297 4199
rect 51859 4168 53297 4196
rect 51859 4165 51871 4168
rect 51813 4159 51871 4165
rect 53285 4165 53297 4168
rect 53331 4196 53343 4199
rect 54941 4199 54999 4205
rect 54941 4196 54953 4199
rect 53331 4168 54953 4196
rect 53331 4165 53343 4168
rect 53285 4159 53343 4165
rect 54941 4165 54953 4168
rect 54987 4196 54999 4199
rect 56413 4199 56471 4205
rect 56413 4196 56425 4199
rect 54987 4168 56425 4196
rect 54987 4165 54999 4168
rect 54941 4159 54999 4165
rect 56413 4165 56425 4168
rect 56459 4196 56471 4199
rect 58161 4199 58219 4205
rect 58161 4196 58173 4199
rect 56459 4168 58173 4196
rect 56459 4165 56471 4168
rect 56413 4159 56471 4165
rect 58161 4165 58173 4168
rect 58207 4196 58219 4199
rect 59449 4199 59507 4205
rect 59449 4196 59461 4199
rect 58207 4168 59461 4196
rect 58207 4165 58219 4168
rect 58161 4159 58219 4165
rect 59449 4165 59461 4168
rect 59495 4196 59507 4199
rect 60918 4196 60924 4208
rect 59495 4168 60924 4196
rect 59495 4165 59507 4168
rect 59449 4159 59507 4165
rect 60918 4156 60924 4168
rect 60976 4196 60982 4208
rect 62393 4199 62451 4205
rect 62393 4196 62405 4199
rect 60976 4168 62405 4196
rect 60976 4156 60982 4168
rect 62393 4165 62405 4168
rect 62439 4196 62451 4199
rect 63865 4199 63923 4205
rect 63865 4196 63877 4199
rect 62439 4168 63877 4196
rect 62439 4165 62451 4168
rect 62393 4159 62451 4165
rect 63865 4165 63877 4168
rect 63911 4165 63923 4199
rect 63865 4159 63923 4165
rect 63954 4156 63960 4208
rect 64012 4205 64018 4208
rect 64012 4199 64040 4205
rect 64028 4165 64040 4199
rect 64012 4159 64040 4165
rect 64012 4156 64018 4159
rect 65334 4156 65340 4208
rect 65392 4196 65398 4208
rect 65392 4168 66484 4196
rect 65392 4156 65398 4168
rect 40681 4131 40739 4137
rect 40681 4097 40693 4131
rect 40727 4097 40739 4131
rect 40681 4091 40739 4097
rect 40862 4088 40868 4140
rect 40920 4128 40926 4140
rect 45370 4128 45376 4140
rect 40920 4100 45376 4128
rect 40920 4088 40926 4100
rect 45370 4088 45376 4100
rect 45428 4088 45434 4140
rect 46566 4088 46572 4140
rect 46624 4128 46630 4140
rect 47146 4131 47204 4137
rect 47146 4128 47158 4131
rect 46624 4100 47158 4128
rect 46624 4088 46630 4100
rect 47146 4097 47158 4100
rect 47192 4097 47204 4131
rect 48225 4131 48283 4137
rect 48225 4128 48237 4131
rect 47146 4091 47204 4097
rect 47320 4100 48237 4128
rect 40770 4060 40776 4072
rect 40604 4032 40776 4060
rect 40770 4020 40776 4032
rect 40828 4020 40834 4072
rect 42334 4060 42340 4072
rect 40880 4032 42340 4060
rect 35434 3992 35440 4004
rect 35176 3964 35440 3992
rect 27522 3884 27528 3936
rect 27580 3884 27586 3936
rect 28626 3884 28632 3936
rect 28684 3884 28690 3936
rect 31018 3884 31024 3936
rect 31076 3884 31082 3936
rect 31110 3884 31116 3936
rect 31168 3924 31174 3936
rect 31662 3924 31668 3936
rect 31168 3896 31668 3924
rect 31168 3884 31174 3896
rect 31662 3884 31668 3896
rect 31720 3884 31726 3936
rect 31849 3927 31907 3933
rect 31849 3893 31861 3927
rect 31895 3924 31907 3927
rect 32214 3924 32220 3936
rect 31895 3896 32220 3924
rect 31895 3893 31907 3896
rect 31849 3887 31907 3893
rect 32214 3884 32220 3896
rect 32272 3884 32278 3936
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 32692 3924 32720 3964
rect 35434 3952 35440 3964
rect 35492 3952 35498 4004
rect 35526 3952 35532 4004
rect 35584 3992 35590 4004
rect 35805 3995 35863 4001
rect 35805 3992 35817 3995
rect 35584 3964 35817 3992
rect 35584 3952 35590 3964
rect 35805 3961 35817 3964
rect 35851 3961 35863 3995
rect 35805 3955 35863 3961
rect 36446 3952 36452 4004
rect 36504 3992 36510 4004
rect 40880 3992 40908 4032
rect 42334 4020 42340 4032
rect 42392 4020 42398 4072
rect 42518 4020 42524 4072
rect 42576 4060 42582 4072
rect 46661 4063 46719 4069
rect 46661 4060 46673 4063
rect 42576 4032 46673 4060
rect 42576 4020 42582 4032
rect 46661 4029 46673 4032
rect 46707 4029 46719 4063
rect 47320 4060 47348 4100
rect 48225 4097 48237 4100
rect 48271 4128 48283 4131
rect 49789 4131 49847 4137
rect 48271 4100 48912 4128
rect 48271 4097 48283 4100
rect 48225 4091 48283 4097
rect 48710 4063 48768 4069
rect 48710 4060 48722 4063
rect 46661 4023 46719 4029
rect 47228 4032 47348 4060
rect 36504 3964 40908 3992
rect 36504 3952 36510 3964
rect 40954 3952 40960 4004
rect 41012 3992 41018 4004
rect 46290 3992 46296 4004
rect 41012 3964 46296 3992
rect 41012 3952 41018 3964
rect 46290 3952 46296 3964
rect 46348 3952 46354 4004
rect 46566 3952 46572 4004
rect 46624 3952 46630 4004
rect 46676 3992 46704 4023
rect 47228 3992 47256 4032
rect 48700 4029 48722 4060
rect 48756 4029 48768 4063
rect 48884 4060 48912 4100
rect 49789 4097 49801 4131
rect 49835 4128 49847 4131
rect 50338 4128 50344 4140
rect 50396 4137 50402 4140
rect 50396 4131 50424 4137
rect 49835 4100 50344 4128
rect 49835 4097 49847 4100
rect 49789 4091 49847 4097
rect 50338 4088 50344 4100
rect 50412 4097 50424 4131
rect 51445 4131 51503 4137
rect 51445 4128 51457 4131
rect 50396 4091 50424 4097
rect 51046 4100 51457 4128
rect 50396 4088 50402 4091
rect 49881 4063 49939 4069
rect 49881 4060 49893 4063
rect 48884 4032 49893 4060
rect 48700 4023 48768 4029
rect 49881 4029 49893 4032
rect 49927 4060 49939 4063
rect 51046 4060 51074 4100
rect 51445 4097 51457 4100
rect 51491 4128 51503 4131
rect 52917 4131 52975 4137
rect 52917 4128 52929 4131
rect 51491 4100 52929 4128
rect 51491 4097 51503 4100
rect 51445 4091 51503 4097
rect 52917 4097 52929 4100
rect 52963 4128 52975 4131
rect 54573 4131 54631 4137
rect 54573 4128 54585 4131
rect 52963 4100 54585 4128
rect 52963 4097 52975 4100
rect 52917 4091 52975 4097
rect 54573 4097 54585 4100
rect 54619 4128 54631 4131
rect 56045 4131 56103 4137
rect 56045 4128 56057 4131
rect 54619 4100 56057 4128
rect 54619 4097 54631 4100
rect 54573 4091 54631 4097
rect 56045 4097 56057 4100
rect 56091 4128 56103 4131
rect 57793 4131 57851 4137
rect 57793 4128 57805 4131
rect 56091 4100 57805 4128
rect 56091 4097 56103 4100
rect 56045 4091 56103 4097
rect 57793 4097 57805 4100
rect 57839 4128 57851 4131
rect 59081 4131 59139 4137
rect 59081 4128 59093 4131
rect 57839 4100 59093 4128
rect 57839 4097 57851 4100
rect 57793 4091 57851 4097
rect 59081 4097 59093 4100
rect 59127 4128 59139 4131
rect 60642 4128 60648 4140
rect 59127 4100 60648 4128
rect 59127 4097 59139 4100
rect 59081 4091 59139 4097
rect 60642 4088 60648 4100
rect 60700 4128 60706 4140
rect 62025 4131 62083 4137
rect 62025 4128 62037 4131
rect 60700 4100 62037 4128
rect 60700 4088 60706 4100
rect 62025 4097 62037 4100
rect 62071 4128 62083 4131
rect 63497 4131 63555 4137
rect 63497 4128 63509 4131
rect 62071 4100 63509 4128
rect 62071 4097 62083 4100
rect 62025 4091 62083 4097
rect 63497 4097 63509 4100
rect 63543 4097 63555 4131
rect 63497 4091 63555 4097
rect 65058 4088 65064 4140
rect 65116 4128 65122 4140
rect 65454 4131 65512 4137
rect 65454 4128 65466 4131
rect 65116 4100 65466 4128
rect 65116 4088 65122 4100
rect 65454 4097 65466 4100
rect 65500 4097 65512 4131
rect 66456 4128 66484 4168
rect 66530 4156 66536 4208
rect 66588 4196 66594 4208
rect 66926 4199 66984 4205
rect 66926 4196 66938 4199
rect 66588 4168 66938 4196
rect 66588 4156 66594 4168
rect 66926 4165 66938 4168
rect 66972 4165 66984 4199
rect 68465 4199 68523 4205
rect 68465 4196 68477 4199
rect 66926 4159 66984 4165
rect 67100 4168 68477 4196
rect 66809 4131 66867 4137
rect 66809 4128 66821 4131
rect 66456 4100 66821 4128
rect 65454 4091 65512 4097
rect 66809 4097 66821 4100
rect 66855 4128 66867 4131
rect 67100 4128 67128 4168
rect 68465 4165 68477 4168
rect 68511 4196 68523 4199
rect 68511 4168 69152 4196
rect 68511 4165 68523 4168
rect 68465 4159 68523 4165
rect 66855 4100 67128 4128
rect 66855 4097 66867 4100
rect 66809 4091 66867 4097
rect 67910 4088 67916 4140
rect 67968 4128 67974 4140
rect 68582 4131 68640 4137
rect 68582 4128 68594 4131
rect 67968 4100 68594 4128
rect 67968 4088 67974 4100
rect 68582 4097 68594 4100
rect 68628 4097 68640 4131
rect 69124 4128 69152 4168
rect 69198 4156 69204 4208
rect 69256 4196 69262 4208
rect 69686 4199 69744 4205
rect 69686 4196 69698 4199
rect 69256 4168 69698 4196
rect 69256 4156 69262 4168
rect 69686 4165 69698 4168
rect 69732 4165 69744 4199
rect 69686 4159 69744 4165
rect 69569 4131 69627 4137
rect 69569 4128 69581 4131
rect 69124 4100 69581 4128
rect 68582 4091 68640 4097
rect 69569 4097 69581 4100
rect 69615 4097 69627 4131
rect 69569 4091 69627 4097
rect 49927 4032 51074 4060
rect 51353 4063 51411 4069
rect 49927 4029 49939 4032
rect 49881 4023 49939 4029
rect 51353 4029 51365 4063
rect 51399 4060 51411 4063
rect 51930 4063 51988 4069
rect 51930 4060 51942 4063
rect 51399 4032 51942 4060
rect 51399 4029 51411 4032
rect 51353 4023 51411 4029
rect 51920 4029 51942 4032
rect 51976 4029 51988 4063
rect 51920 4023 51988 4029
rect 46676 3964 47256 3992
rect 47305 3995 47363 4001
rect 47305 3961 47317 3995
rect 47351 3992 47363 3995
rect 48590 3992 48596 4004
rect 47351 3964 48596 3992
rect 47351 3961 47363 3964
rect 47305 3955 47363 3961
rect 48590 3952 48596 3964
rect 48648 3952 48654 4004
rect 32456 3896 32720 3924
rect 32769 3927 32827 3933
rect 32456 3884 32462 3896
rect 32769 3893 32781 3927
rect 32815 3924 32827 3927
rect 33134 3924 33140 3936
rect 32815 3896 33140 3924
rect 32815 3893 32827 3896
rect 32769 3887 32827 3893
rect 33134 3884 33140 3896
rect 33192 3884 33198 3936
rect 33413 3927 33471 3933
rect 33413 3893 33425 3927
rect 33459 3924 33471 3927
rect 33502 3924 33508 3936
rect 33459 3896 33508 3924
rect 33459 3893 33471 3896
rect 33413 3887 33471 3893
rect 33502 3884 33508 3896
rect 33560 3884 33566 3936
rect 33778 3884 33784 3936
rect 33836 3924 33842 3936
rect 34054 3924 34060 3936
rect 33836 3896 34060 3924
rect 33836 3884 33842 3896
rect 34054 3884 34060 3896
rect 34112 3884 34118 3936
rect 36170 3884 36176 3936
rect 36228 3924 36234 3936
rect 47578 3924 47584 3936
rect 36228 3896 47584 3924
rect 36228 3884 36234 3896
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 48130 3884 48136 3936
rect 48188 3924 48194 3936
rect 48700 3924 48728 4023
rect 48869 3995 48927 4001
rect 48869 3961 48881 3995
rect 48915 3992 48927 3995
rect 50525 3995 50583 4001
rect 48915 3964 50016 3992
rect 48915 3961 48927 3964
rect 48869 3955 48927 3961
rect 48188 3896 48728 3924
rect 49988 3924 50016 3964
rect 50525 3961 50537 3995
rect 50571 3992 50583 3995
rect 51074 3992 51080 4004
rect 50571 3964 51080 3992
rect 50571 3961 50583 3964
rect 50525 3955 50583 3961
rect 51074 3952 51080 3964
rect 51132 3952 51138 4004
rect 51442 3992 51448 4004
rect 51184 3964 51448 3992
rect 51184 3924 51212 3964
rect 51442 3952 51448 3964
rect 51500 3952 51506 4004
rect 49988 3896 51212 3924
rect 51920 3924 51948 4023
rect 53374 4020 53380 4072
rect 53432 4069 53438 4072
rect 53432 4063 53460 4069
rect 53448 4029 53460 4063
rect 53432 4023 53460 4029
rect 54481 4063 54539 4069
rect 54481 4029 54493 4063
rect 54527 4060 54539 4063
rect 55030 4060 55036 4072
rect 55088 4069 55094 4072
rect 55088 4063 55116 4069
rect 54527 4032 55036 4060
rect 54527 4029 54539 4032
rect 54481 4023 54539 4029
rect 53432 4020 53438 4023
rect 55030 4020 55036 4032
rect 55104 4029 55116 4063
rect 55088 4023 55116 4029
rect 55953 4063 56011 4069
rect 55953 4029 55965 4063
rect 55999 4060 56011 4063
rect 56502 4060 56508 4072
rect 56560 4069 56566 4072
rect 56560 4063 56588 4069
rect 55999 4032 56508 4060
rect 55999 4029 56011 4032
rect 55953 4023 56011 4029
rect 55088 4020 55094 4023
rect 56502 4020 56508 4032
rect 56576 4029 56588 4063
rect 56560 4023 56588 4029
rect 56560 4020 56566 4023
rect 58250 4020 58256 4072
rect 58308 4069 58314 4072
rect 58308 4063 58336 4069
rect 58324 4029 58336 4063
rect 58308 4023 58336 4029
rect 58308 4020 58314 4023
rect 59170 4020 59176 4072
rect 59228 4060 59234 4072
rect 59566 4063 59624 4069
rect 59566 4060 59578 4063
rect 59228 4032 59578 4060
rect 59228 4020 59234 4032
rect 59566 4029 59578 4032
rect 59612 4029 59624 4063
rect 59566 4023 59624 4029
rect 62298 4020 62304 4072
rect 62356 4060 62362 4072
rect 62510 4063 62568 4069
rect 62510 4060 62522 4063
rect 62356 4032 62522 4060
rect 62356 4020 62362 4032
rect 62510 4029 62522 4032
rect 62556 4029 62568 4063
rect 62510 4023 62568 4029
rect 64969 4063 65027 4069
rect 64969 4029 64981 4063
rect 65015 4060 65027 4063
rect 66441 4063 66499 4069
rect 66441 4060 66453 4063
rect 65015 4032 66453 4060
rect 65015 4029 65027 4032
rect 64969 4023 65027 4029
rect 66441 4029 66453 4032
rect 66487 4060 66499 4063
rect 68097 4063 68155 4069
rect 68097 4060 68109 4063
rect 66487 4032 68109 4060
rect 66487 4029 66499 4032
rect 66441 4023 66499 4029
rect 68097 4029 68109 4032
rect 68143 4060 68155 4063
rect 69201 4063 69259 4069
rect 69201 4060 69213 4063
rect 68143 4032 69213 4060
rect 68143 4029 68155 4032
rect 68097 4023 68155 4029
rect 69201 4029 69213 4032
rect 69247 4029 69259 4063
rect 69201 4023 69259 4029
rect 52089 3995 52147 4001
rect 52089 3961 52101 3995
rect 52135 3992 52147 3995
rect 55217 3995 55275 4001
rect 52135 3964 54892 3992
rect 52135 3961 52147 3964
rect 52089 3955 52147 3961
rect 54864 3936 54892 3964
rect 55217 3961 55229 3995
rect 55263 3992 55275 3995
rect 57422 3992 57428 4004
rect 55263 3964 57428 3992
rect 55263 3961 55275 3964
rect 55217 3955 55275 3961
rect 57422 3952 57428 3964
rect 57480 3952 57486 4004
rect 59725 3995 59783 4001
rect 59725 3961 59737 3995
rect 59771 3992 59783 3995
rect 61654 3992 61660 4004
rect 59771 3964 61660 3992
rect 59771 3961 59783 3964
rect 59725 3955 59783 3961
rect 61654 3952 61660 3964
rect 61712 3952 61718 4004
rect 63862 3952 63868 4004
rect 63920 3992 63926 4004
rect 64984 3992 65012 4023
rect 63920 3964 65012 3992
rect 68741 3995 68799 4001
rect 63920 3952 63926 3964
rect 68741 3961 68753 3995
rect 68787 3992 68799 3995
rect 70578 3992 70584 4004
rect 68787 3964 70584 3992
rect 68787 3961 68799 3964
rect 68741 3955 68799 3961
rect 70578 3952 70584 3964
rect 70636 3952 70642 4004
rect 52362 3924 52368 3936
rect 51920 3896 52368 3924
rect 48188 3884 48194 3896
rect 52362 3884 52368 3896
rect 52420 3884 52426 3936
rect 53561 3927 53619 3933
rect 53561 3893 53573 3927
rect 53607 3924 53619 3927
rect 54018 3924 54024 3936
rect 53607 3896 54024 3924
rect 53607 3893 53619 3896
rect 53561 3887 53619 3893
rect 54018 3884 54024 3896
rect 54076 3884 54082 3936
rect 54846 3884 54852 3936
rect 54904 3884 54910 3936
rect 56689 3927 56747 3933
rect 56689 3893 56701 3927
rect 56735 3924 56747 3927
rect 57606 3924 57612 3936
rect 56735 3896 57612 3924
rect 56735 3893 56747 3896
rect 56689 3887 56747 3893
rect 57606 3884 57612 3896
rect 57664 3884 57670 3936
rect 58434 3884 58440 3936
rect 58492 3884 58498 3936
rect 62666 3884 62672 3936
rect 62724 3884 62730 3936
rect 64141 3927 64199 3933
rect 64141 3893 64153 3927
rect 64187 3924 64199 3927
rect 65334 3924 65340 3936
rect 64187 3896 65340 3924
rect 64187 3893 64199 3896
rect 64141 3887 64199 3893
rect 65334 3884 65340 3896
rect 65392 3884 65398 3936
rect 65613 3927 65671 3933
rect 65613 3893 65625 3927
rect 65659 3924 65671 3927
rect 66990 3924 66996 3936
rect 65659 3896 66996 3924
rect 65659 3893 65671 3896
rect 65613 3887 65671 3893
rect 66990 3884 66996 3896
rect 67048 3884 67054 3936
rect 67085 3927 67143 3933
rect 67085 3893 67097 3927
rect 67131 3924 67143 3927
rect 69382 3924 69388 3936
rect 67131 3896 69388 3924
rect 67131 3893 67143 3896
rect 67085 3887 67143 3893
rect 69382 3884 69388 3896
rect 69440 3884 69446 3936
rect 69845 3927 69903 3933
rect 69845 3893 69857 3927
rect 69891 3924 69903 3927
rect 71406 3924 71412 3936
rect 69891 3896 71412 3924
rect 69891 3893 69903 3896
rect 69845 3887 69903 3893
rect 71406 3884 71412 3896
rect 71464 3884 71470 3936
rect 1012 3834 74980 3856
rect 1012 3782 1858 3834
rect 1910 3782 1922 3834
rect 1974 3782 1986 3834
rect 2038 3782 2050 3834
rect 2102 3782 2114 3834
rect 2166 3782 11858 3834
rect 11910 3782 11922 3834
rect 11974 3782 11986 3834
rect 12038 3782 12050 3834
rect 12102 3782 12114 3834
rect 12166 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 21986 3834
rect 22038 3782 22050 3834
rect 22102 3782 22114 3834
rect 22166 3782 31858 3834
rect 31910 3782 31922 3834
rect 31974 3782 31986 3834
rect 32038 3782 32050 3834
rect 32102 3782 32114 3834
rect 32166 3782 41858 3834
rect 41910 3782 41922 3834
rect 41974 3782 41986 3834
rect 42038 3782 42050 3834
rect 42102 3782 42114 3834
rect 42166 3782 51858 3834
rect 51910 3782 51922 3834
rect 51974 3782 51986 3834
rect 52038 3782 52050 3834
rect 52102 3782 52114 3834
rect 52166 3782 61858 3834
rect 61910 3782 61922 3834
rect 61974 3782 61986 3834
rect 62038 3782 62050 3834
rect 62102 3782 62114 3834
rect 62166 3782 71858 3834
rect 71910 3782 71922 3834
rect 71974 3782 71986 3834
rect 72038 3782 72050 3834
rect 72102 3782 72114 3834
rect 72166 3782 74980 3834
rect 1012 3760 74980 3782
rect 32306 3720 32312 3732
rect 31312 3692 32312 3720
rect 26878 3544 26884 3596
rect 26936 3544 26942 3596
rect 28629 3587 28687 3593
rect 28629 3584 28641 3587
rect 27080 3556 28641 3584
rect 27080 3525 27108 3556
rect 28629 3553 28641 3556
rect 28675 3553 28687 3587
rect 28629 3547 28687 3553
rect 29914 3544 29920 3596
rect 29972 3584 29978 3596
rect 30469 3587 30527 3593
rect 30469 3584 30481 3587
rect 29972 3556 30481 3584
rect 29972 3544 29978 3556
rect 30469 3553 30481 3556
rect 30515 3584 30527 3587
rect 30650 3584 30656 3596
rect 30515 3556 30656 3584
rect 30515 3553 30527 3556
rect 30469 3547 30527 3553
rect 30650 3544 30656 3556
rect 30708 3584 30714 3596
rect 31312 3593 31340 3692
rect 31687 3661 31693 3664
rect 31665 3655 31693 3661
rect 31665 3621 31677 3655
rect 31665 3615 31693 3621
rect 31687 3612 31693 3615
rect 31745 3612 31751 3664
rect 31297 3587 31355 3593
rect 31297 3584 31309 3587
rect 30708 3556 31309 3584
rect 30708 3544 30714 3556
rect 31297 3553 31309 3556
rect 31343 3553 31355 3587
rect 31297 3547 31355 3553
rect 31386 3544 31392 3596
rect 31444 3544 31450 3596
rect 31478 3544 31484 3596
rect 31536 3593 31542 3596
rect 32048 3593 32076 3692
rect 32306 3680 32312 3692
rect 32364 3680 32370 3732
rect 32769 3723 32827 3729
rect 32769 3689 32781 3723
rect 32815 3720 32827 3723
rect 33318 3720 33324 3732
rect 32815 3692 33324 3720
rect 32815 3689 32827 3692
rect 32769 3683 32827 3689
rect 33318 3680 33324 3692
rect 33376 3680 33382 3732
rect 34425 3723 34483 3729
rect 34425 3689 34437 3723
rect 34471 3720 34483 3723
rect 34790 3720 34796 3732
rect 34471 3692 34796 3720
rect 34471 3689 34483 3692
rect 34425 3683 34483 3689
rect 34790 3680 34796 3692
rect 34848 3720 34854 3732
rect 35713 3723 35771 3729
rect 35713 3720 35725 3723
rect 34848 3692 35725 3720
rect 34848 3680 34854 3692
rect 35713 3689 35725 3692
rect 35759 3720 35771 3723
rect 35986 3720 35992 3732
rect 35759 3692 35992 3720
rect 35759 3689 35771 3692
rect 35713 3683 35771 3689
rect 35986 3680 35992 3692
rect 36044 3680 36050 3732
rect 37921 3723 37979 3729
rect 37921 3689 37933 3723
rect 37967 3720 37979 3723
rect 40862 3720 40868 3732
rect 37967 3692 40868 3720
rect 37967 3689 37979 3692
rect 37921 3683 37979 3689
rect 40862 3680 40868 3692
rect 40920 3680 40926 3732
rect 41322 3680 41328 3732
rect 41380 3720 41386 3732
rect 60642 3720 60648 3732
rect 41380 3692 60648 3720
rect 41380 3680 41386 3692
rect 60642 3680 60648 3692
rect 60700 3680 60706 3732
rect 64782 3720 64788 3732
rect 61672 3692 64788 3720
rect 32398 3612 32404 3664
rect 32456 3612 32462 3664
rect 32950 3652 32956 3664
rect 32876 3624 32956 3652
rect 32876 3593 32904 3624
rect 32950 3612 32956 3624
rect 33008 3652 33014 3664
rect 33962 3652 33968 3664
rect 33008 3624 33968 3652
rect 33008 3612 33014 3624
rect 33962 3612 33968 3624
rect 34020 3612 34026 3664
rect 34701 3655 34759 3661
rect 34701 3652 34713 3655
rect 34348 3624 34713 3652
rect 31536 3587 31564 3593
rect 31552 3553 31564 3587
rect 31536 3547 31564 3553
rect 32033 3587 32091 3593
rect 32033 3553 32045 3587
rect 32079 3584 32091 3587
rect 32861 3587 32919 3593
rect 32079 3556 32720 3584
rect 32079 3553 32091 3556
rect 32033 3547 32091 3553
rect 31536 3544 31542 3547
rect 27065 3519 27123 3525
rect 27065 3485 27077 3519
rect 27111 3485 27123 3519
rect 27065 3479 27123 3485
rect 27154 3476 27160 3528
rect 27212 3476 27218 3528
rect 27982 3476 27988 3528
rect 28040 3476 28046 3528
rect 29181 3519 29239 3525
rect 29181 3516 29193 3519
rect 28092 3488 29193 3516
rect 26602 3408 26608 3460
rect 26660 3448 26666 3460
rect 28092 3448 28120 3488
rect 29181 3485 29193 3488
rect 29227 3485 29239 3519
rect 29181 3479 29239 3485
rect 29457 3519 29515 3525
rect 29457 3485 29469 3519
rect 29503 3485 29515 3519
rect 29457 3479 29515 3485
rect 30193 3519 30251 3525
rect 30193 3485 30205 3519
rect 30239 3516 30251 3519
rect 31021 3519 31079 3525
rect 31021 3516 31033 3519
rect 30239 3488 31033 3516
rect 30239 3485 30251 3488
rect 30193 3479 30251 3485
rect 31021 3485 31033 3488
rect 31067 3516 31079 3519
rect 31757 3519 31815 3525
rect 31757 3516 31769 3519
rect 31067 3488 31769 3516
rect 31067 3485 31079 3488
rect 31021 3479 31079 3485
rect 31757 3485 31769 3488
rect 31803 3485 31815 3519
rect 31757 3479 31815 3485
rect 32242 3519 32300 3525
rect 32242 3485 32254 3519
rect 32288 3516 32300 3519
rect 32582 3516 32588 3528
rect 32288 3488 32588 3516
rect 32288 3485 32300 3488
rect 32242 3479 32300 3485
rect 26660 3420 28120 3448
rect 28537 3451 28595 3457
rect 26660 3408 26666 3420
rect 28537 3417 28549 3451
rect 28583 3448 28595 3451
rect 29472 3448 29500 3479
rect 28583 3420 29500 3448
rect 28583 3417 28595 3420
rect 28537 3411 28595 3417
rect 29730 3408 29736 3460
rect 29788 3408 29794 3460
rect 30101 3451 30159 3457
rect 30101 3417 30113 3451
rect 30147 3448 30159 3451
rect 30282 3448 30288 3460
rect 30147 3420 30288 3448
rect 30147 3417 30159 3420
rect 30101 3411 30159 3417
rect 30282 3408 30288 3420
rect 30340 3448 30346 3460
rect 30653 3451 30711 3457
rect 30653 3448 30665 3451
rect 30340 3420 30665 3448
rect 30340 3408 30346 3420
rect 30653 3417 30665 3420
rect 30699 3417 30711 3451
rect 30653 3411 30711 3417
rect 30926 3408 30932 3460
rect 30984 3408 30990 3460
rect 31772 3448 31800 3479
rect 32582 3476 32588 3488
rect 32640 3476 32646 3528
rect 32692 3516 32720 3556
rect 32861 3553 32873 3587
rect 32907 3553 32919 3587
rect 32861 3547 32919 3553
rect 33042 3544 33048 3596
rect 33100 3584 33106 3596
rect 33100 3556 34100 3584
rect 33100 3544 33106 3556
rect 33137 3519 33195 3525
rect 33137 3516 33149 3519
rect 32692 3488 33149 3516
rect 33137 3485 33149 3488
rect 33183 3485 33195 3519
rect 33137 3479 33195 3485
rect 33318 3476 33324 3528
rect 33376 3525 33382 3528
rect 33376 3519 33404 3525
rect 33392 3485 33404 3519
rect 33376 3479 33404 3485
rect 33597 3519 33655 3525
rect 33597 3485 33609 3519
rect 33643 3516 33655 3519
rect 33962 3516 33968 3528
rect 33643 3488 33968 3516
rect 33643 3485 33655 3488
rect 33597 3479 33655 3485
rect 33376 3476 33382 3479
rect 33962 3476 33968 3488
rect 34020 3476 34026 3528
rect 34072 3516 34100 3556
rect 34348 3516 34376 3624
rect 34701 3621 34713 3624
rect 34747 3621 34759 3655
rect 35529 3655 35587 3661
rect 35529 3652 35541 3655
rect 34701 3615 34759 3621
rect 34875 3624 35541 3652
rect 34875 3593 34903 3624
rect 35529 3621 35541 3624
rect 35575 3652 35587 3655
rect 36078 3652 36084 3664
rect 35575 3624 36084 3652
rect 35575 3621 35587 3624
rect 35529 3615 35587 3621
rect 36078 3612 36084 3624
rect 36136 3612 36142 3664
rect 36188 3624 45692 3652
rect 34860 3587 34918 3593
rect 34860 3553 34872 3587
rect 34906 3553 34918 3587
rect 34860 3547 34918 3553
rect 35250 3544 35256 3596
rect 35308 3584 35314 3596
rect 36188 3593 36216 3624
rect 35345 3587 35403 3593
rect 35345 3584 35357 3587
rect 35308 3556 35357 3584
rect 35308 3544 35314 3556
rect 35345 3553 35357 3556
rect 35391 3553 35403 3587
rect 35345 3547 35403 3553
rect 36173 3587 36231 3593
rect 36173 3553 36185 3587
rect 36219 3553 36231 3587
rect 40126 3584 40132 3596
rect 36173 3547 36231 3553
rect 36280 3556 40132 3584
rect 34072 3488 34376 3516
rect 35069 3519 35127 3525
rect 35069 3485 35081 3519
rect 35115 3485 35127 3519
rect 35069 3479 35127 3485
rect 32950 3448 32956 3460
rect 31772 3420 32956 3448
rect 32950 3408 32956 3420
rect 33008 3408 33014 3460
rect 33244 3420 34008 3448
rect 27798 3340 27804 3392
rect 27856 3340 27862 3392
rect 30561 3383 30619 3389
rect 30561 3349 30573 3383
rect 30607 3380 30619 3383
rect 31386 3380 31392 3392
rect 30607 3352 31392 3380
rect 30607 3349 30619 3352
rect 30561 3343 30619 3349
rect 31386 3340 31392 3352
rect 31444 3380 31450 3392
rect 33244 3389 33272 3420
rect 33980 3392 34008 3420
rect 34054 3408 34060 3460
rect 34112 3457 34118 3460
rect 34112 3451 34140 3457
rect 34128 3417 34140 3451
rect 35084 3448 35112 3479
rect 35342 3448 35348 3460
rect 35084 3420 35348 3448
rect 34112 3411 34140 3417
rect 34112 3408 34118 3411
rect 35342 3408 35348 3420
rect 35400 3408 35406 3460
rect 35434 3408 35440 3460
rect 35492 3448 35498 3460
rect 36280 3448 36308 3556
rect 40126 3544 40132 3556
rect 40184 3544 40190 3596
rect 41325 3587 41383 3593
rect 40236 3556 40448 3584
rect 36354 3476 36360 3528
rect 36412 3476 36418 3528
rect 36909 3519 36967 3525
rect 36909 3485 36921 3519
rect 36955 3516 36967 3519
rect 40236 3516 40264 3556
rect 36955 3488 40264 3516
rect 40420 3516 40448 3556
rect 41325 3553 41337 3587
rect 41371 3584 41383 3587
rect 45664 3584 45692 3624
rect 46566 3612 46572 3664
rect 46624 3652 46630 3664
rect 46753 3655 46811 3661
rect 46753 3652 46765 3655
rect 46624 3624 46765 3652
rect 46624 3612 46630 3624
rect 46753 3621 46765 3624
rect 46799 3652 46811 3655
rect 48130 3652 48136 3664
rect 46799 3624 48136 3652
rect 46799 3621 46811 3624
rect 46753 3615 46811 3621
rect 48130 3612 48136 3624
rect 48188 3612 48194 3664
rect 51074 3612 51080 3664
rect 51132 3652 51138 3664
rect 53098 3652 53104 3664
rect 51132 3624 53104 3652
rect 51132 3612 51138 3624
rect 53098 3612 53104 3624
rect 53156 3612 53162 3664
rect 58434 3612 58440 3664
rect 58492 3652 58498 3664
rect 61562 3652 61568 3664
rect 58492 3624 61568 3652
rect 58492 3612 58498 3624
rect 61562 3612 61568 3624
rect 61620 3612 61626 3664
rect 41371 3556 45600 3584
rect 45664 3556 57744 3584
rect 41371 3553 41383 3556
rect 41325 3547 41383 3553
rect 45462 3516 45468 3528
rect 40420 3488 45468 3516
rect 36955 3485 36967 3488
rect 36909 3479 36967 3485
rect 45462 3476 45468 3488
rect 45520 3476 45526 3528
rect 45572 3516 45600 3556
rect 50982 3516 50988 3528
rect 45572 3488 50988 3516
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 51442 3476 51448 3528
rect 51500 3516 51506 3528
rect 52270 3516 52276 3528
rect 51500 3488 52276 3516
rect 51500 3476 51506 3488
rect 52270 3476 52276 3488
rect 52328 3476 52334 3528
rect 57606 3476 57612 3528
rect 57664 3476 57670 3528
rect 57716 3516 57744 3556
rect 57790 3544 57796 3596
rect 57848 3584 57854 3596
rect 61672 3584 61700 3692
rect 64782 3680 64788 3692
rect 64840 3680 64846 3732
rect 64966 3680 64972 3732
rect 65024 3680 65030 3732
rect 66530 3680 66536 3732
rect 66588 3680 66594 3732
rect 67910 3680 67916 3732
rect 67968 3720 67974 3732
rect 68097 3723 68155 3729
rect 68097 3720 68109 3723
rect 67968 3692 68109 3720
rect 67968 3680 67974 3692
rect 68097 3689 68109 3692
rect 68143 3689 68155 3723
rect 68097 3683 68155 3689
rect 69198 3680 69204 3732
rect 69256 3680 69262 3732
rect 62117 3655 62175 3661
rect 62117 3621 62129 3655
rect 62163 3652 62175 3655
rect 62298 3652 62304 3664
rect 62163 3624 62304 3652
rect 62163 3621 62175 3624
rect 62117 3615 62175 3621
rect 62298 3612 62304 3624
rect 62356 3612 62362 3664
rect 63494 3612 63500 3664
rect 63552 3652 63558 3664
rect 63589 3655 63647 3661
rect 63589 3652 63601 3655
rect 63552 3624 63601 3652
rect 63552 3612 63558 3624
rect 63589 3621 63601 3624
rect 63635 3652 63647 3655
rect 63954 3652 63960 3664
rect 63635 3624 63960 3652
rect 63635 3621 63647 3624
rect 63589 3615 63647 3621
rect 63954 3612 63960 3624
rect 64012 3612 64018 3664
rect 65705 3655 65763 3661
rect 65705 3621 65717 3655
rect 65751 3652 65763 3655
rect 66898 3652 66904 3664
rect 65751 3624 66904 3652
rect 65751 3621 65763 3624
rect 65705 3615 65763 3621
rect 66898 3612 66904 3624
rect 66956 3612 66962 3664
rect 57848 3556 61700 3584
rect 64325 3587 64383 3593
rect 57848 3544 57854 3556
rect 64325 3553 64337 3587
rect 64371 3584 64383 3587
rect 67542 3584 67548 3596
rect 64371 3556 67548 3584
rect 64371 3553 64383 3556
rect 64325 3547 64383 3553
rect 67542 3544 67548 3556
rect 67600 3544 67606 3596
rect 61470 3516 61476 3528
rect 57716 3488 61476 3516
rect 61470 3476 61476 3488
rect 61528 3476 61534 3528
rect 63773 3519 63831 3525
rect 63773 3485 63785 3519
rect 63819 3516 63831 3519
rect 65426 3516 65432 3528
rect 63819 3488 65432 3516
rect 63819 3485 63831 3488
rect 63773 3479 63831 3485
rect 65426 3476 65432 3488
rect 65484 3476 65490 3528
rect 35492 3420 36308 3448
rect 35492 3408 35498 3420
rect 36538 3408 36544 3460
rect 36596 3408 36602 3460
rect 38013 3451 38071 3457
rect 38013 3417 38025 3451
rect 38059 3448 38071 3451
rect 38378 3448 38384 3460
rect 38059 3420 38384 3448
rect 38059 3417 38071 3420
rect 38013 3411 38071 3417
rect 38378 3408 38384 3420
rect 38436 3408 38442 3460
rect 40218 3448 40224 3460
rect 38764 3420 40224 3448
rect 32125 3383 32183 3389
rect 32125 3380 32137 3383
rect 31444 3352 32137 3380
rect 31444 3340 31450 3352
rect 32125 3349 32137 3352
rect 32171 3380 32183 3383
rect 33229 3383 33287 3389
rect 33229 3380 33241 3383
rect 32171 3352 33241 3380
rect 32171 3349 32183 3352
rect 32125 3343 32183 3349
rect 33229 3349 33241 3352
rect 33275 3349 33287 3383
rect 33229 3343 33287 3349
rect 33410 3340 33416 3392
rect 33468 3380 33474 3392
rect 33505 3383 33563 3389
rect 33505 3380 33517 3383
rect 33468 3352 33517 3380
rect 33468 3340 33474 3352
rect 33505 3349 33517 3352
rect 33551 3349 33563 3383
rect 33505 3343 33563 3349
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 33873 3383 33931 3389
rect 33873 3380 33885 3383
rect 33652 3352 33885 3380
rect 33652 3340 33658 3352
rect 33873 3349 33885 3352
rect 33919 3349 33931 3383
rect 33873 3343 33931 3349
rect 33962 3340 33968 3392
rect 34020 3340 34026 3392
rect 34241 3383 34299 3389
rect 34241 3349 34253 3383
rect 34287 3380 34299 3383
rect 34606 3380 34612 3392
rect 34287 3352 34612 3380
rect 34287 3349 34299 3352
rect 34241 3343 34299 3349
rect 34606 3340 34612 3352
rect 34664 3340 34670 3392
rect 34974 3340 34980 3392
rect 35032 3340 35038 3392
rect 35066 3340 35072 3392
rect 35124 3380 35130 3392
rect 35526 3380 35532 3392
rect 35124 3352 35532 3380
rect 35124 3340 35130 3352
rect 35526 3340 35532 3352
rect 35584 3340 35590 3392
rect 35710 3340 35716 3392
rect 35768 3380 35774 3392
rect 38764 3380 38792 3420
rect 40218 3408 40224 3420
rect 40276 3408 40282 3460
rect 40310 3408 40316 3460
rect 40368 3448 40374 3460
rect 41506 3448 41512 3460
rect 40368 3420 41512 3448
rect 40368 3408 40374 3420
rect 41506 3408 41512 3420
rect 41564 3408 41570 3460
rect 41598 3408 41604 3460
rect 41656 3408 41662 3460
rect 42242 3408 42248 3460
rect 42300 3448 42306 3460
rect 42300 3420 46244 3448
rect 42300 3408 42306 3420
rect 35768 3352 38792 3380
rect 35768 3340 35774 3352
rect 38838 3340 38844 3392
rect 38896 3380 38902 3392
rect 46106 3380 46112 3392
rect 38896 3352 46112 3380
rect 38896 3340 38902 3352
rect 46106 3340 46112 3352
rect 46164 3340 46170 3392
rect 46216 3380 46244 3420
rect 46290 3408 46296 3460
rect 46348 3448 46354 3460
rect 48038 3448 48044 3460
rect 46348 3420 48044 3448
rect 46348 3408 46354 3420
rect 48038 3408 48044 3420
rect 48096 3408 48102 3460
rect 48130 3408 48136 3460
rect 48188 3448 48194 3460
rect 58710 3448 58716 3460
rect 48188 3420 58716 3448
rect 48188 3408 48194 3420
rect 58710 3408 58716 3420
rect 58768 3408 58774 3460
rect 58805 3451 58863 3457
rect 58805 3417 58817 3451
rect 58851 3448 58863 3451
rect 58894 3448 58900 3460
rect 58851 3420 58900 3448
rect 58851 3417 58863 3420
rect 58805 3411 58863 3417
rect 58894 3408 58900 3420
rect 58952 3408 58958 3460
rect 62574 3448 62580 3460
rect 61948 3420 62580 3448
rect 52730 3380 52736 3392
rect 46216 3352 52736 3380
rect 52730 3340 52736 3352
rect 52788 3340 52794 3392
rect 53006 3340 53012 3392
rect 53064 3340 53070 3392
rect 59170 3340 59176 3392
rect 59228 3340 59234 3392
rect 60550 3340 60556 3392
rect 60608 3340 60614 3392
rect 60642 3340 60648 3392
rect 60700 3380 60706 3392
rect 61948 3380 61976 3420
rect 62574 3408 62580 3420
rect 62632 3408 62638 3460
rect 65886 3408 65892 3460
rect 65944 3408 65950 3460
rect 60700 3352 61976 3380
rect 60700 3340 60706 3352
rect 62390 3340 62396 3392
rect 62448 3380 62454 3392
rect 69106 3380 69112 3392
rect 62448 3352 69112 3380
rect 62448 3340 62454 3352
rect 69106 3340 69112 3352
rect 69164 3340 69170 3392
rect 1012 3290 74980 3312
rect 1012 3238 4210 3290
rect 4262 3238 4274 3290
rect 4326 3238 4338 3290
rect 4390 3238 4402 3290
rect 4454 3238 4466 3290
rect 4518 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 24466 3290
rect 24518 3238 34210 3290
rect 34262 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 44210 3290
rect 44262 3238 44274 3290
rect 44326 3238 44338 3290
rect 44390 3238 44402 3290
rect 44454 3238 44466 3290
rect 44518 3238 54210 3290
rect 54262 3238 54274 3290
rect 54326 3238 54338 3290
rect 54390 3238 54402 3290
rect 54454 3238 54466 3290
rect 54518 3238 64210 3290
rect 64262 3238 64274 3290
rect 64326 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 74210 3290
rect 74262 3238 74274 3290
rect 74326 3238 74338 3290
rect 74390 3238 74402 3290
rect 74454 3238 74466 3290
rect 74518 3238 74980 3290
rect 1012 3216 74980 3238
rect 27982 3136 27988 3188
rect 28040 3176 28046 3188
rect 28077 3179 28135 3185
rect 28077 3176 28089 3179
rect 28040 3148 28089 3176
rect 28040 3136 28046 3148
rect 28077 3145 28089 3148
rect 28123 3145 28135 3179
rect 28077 3139 28135 3145
rect 29454 3136 29460 3188
rect 29512 3176 29518 3188
rect 29549 3179 29607 3185
rect 29549 3176 29561 3179
rect 29512 3148 29561 3176
rect 29512 3136 29518 3148
rect 29549 3145 29561 3148
rect 29595 3145 29607 3179
rect 31294 3176 31300 3188
rect 29549 3139 29607 3145
rect 30944 3148 31300 3176
rect 26421 3111 26479 3117
rect 26421 3077 26433 3111
rect 26467 3108 26479 3111
rect 30944 3108 30972 3148
rect 31294 3136 31300 3148
rect 31352 3136 31358 3188
rect 31849 3179 31907 3185
rect 31849 3145 31861 3179
rect 31895 3176 31907 3179
rect 32582 3176 32588 3188
rect 31895 3148 32588 3176
rect 31895 3145 31907 3148
rect 31849 3139 31907 3145
rect 32582 3136 32588 3148
rect 32640 3136 32646 3188
rect 32766 3136 32772 3188
rect 32824 3136 32830 3188
rect 33137 3179 33195 3185
rect 33137 3145 33149 3179
rect 33183 3176 33195 3179
rect 33686 3176 33692 3188
rect 33183 3148 33692 3176
rect 33183 3145 33195 3148
rect 33137 3139 33195 3145
rect 33686 3136 33692 3148
rect 33744 3136 33750 3188
rect 33778 3136 33784 3188
rect 33836 3176 33842 3188
rect 39758 3176 39764 3188
rect 33836 3148 39764 3176
rect 33836 3136 33842 3148
rect 39758 3136 39764 3148
rect 39816 3136 39822 3188
rect 41969 3179 42027 3185
rect 41969 3145 41981 3179
rect 42015 3176 42027 3179
rect 42242 3176 42248 3188
rect 42015 3148 42248 3176
rect 42015 3145 42027 3148
rect 41969 3139 42027 3145
rect 42242 3136 42248 3148
rect 42300 3136 42306 3188
rect 44545 3179 44603 3185
rect 44545 3145 44557 3179
rect 44591 3176 44603 3179
rect 45002 3176 45008 3188
rect 44591 3148 45008 3176
rect 44591 3145 44603 3148
rect 44545 3139 44603 3145
rect 45002 3136 45008 3148
rect 45060 3136 45066 3188
rect 45373 3179 45431 3185
rect 45373 3145 45385 3179
rect 45419 3176 45431 3179
rect 50890 3176 50896 3188
rect 45419 3148 50896 3176
rect 45419 3145 45431 3148
rect 45373 3139 45431 3145
rect 50890 3136 50896 3148
rect 50948 3136 50954 3188
rect 50982 3136 50988 3188
rect 51040 3176 51046 3188
rect 51718 3176 51724 3188
rect 51040 3148 51724 3176
rect 51040 3136 51046 3148
rect 51718 3136 51724 3148
rect 51776 3136 51782 3188
rect 57790 3176 57796 3188
rect 55140 3148 57796 3176
rect 26467 3080 30972 3108
rect 26467 3077 26479 3080
rect 26421 3071 26479 3077
rect 31018 3068 31024 3120
rect 31076 3108 31082 3120
rect 33318 3108 33324 3120
rect 31076 3080 33324 3108
rect 31076 3068 31082 3080
rect 33318 3068 33324 3080
rect 33376 3068 33382 3120
rect 34054 3068 34060 3120
rect 34112 3068 34118 3120
rect 34701 3111 34759 3117
rect 34701 3077 34713 3111
rect 34747 3108 34759 3111
rect 35526 3108 35532 3120
rect 34747 3080 35532 3108
rect 34747 3077 34759 3080
rect 34701 3071 34759 3077
rect 35526 3068 35532 3080
rect 35584 3068 35590 3120
rect 44910 3108 44916 3120
rect 35728 3080 44916 3108
rect 25682 3000 25688 3052
rect 25740 3000 25746 3052
rect 26694 3000 26700 3052
rect 26752 3000 26758 3052
rect 27433 3043 27491 3049
rect 27433 3009 27445 3043
rect 27479 3040 27491 3043
rect 28626 3040 28632 3052
rect 27479 3012 28632 3040
rect 27479 3009 27491 3012
rect 27433 3003 27491 3009
rect 28626 3000 28632 3012
rect 28684 3000 28690 3052
rect 28721 3043 28779 3049
rect 28721 3009 28733 3043
rect 28767 3040 28779 3043
rect 29914 3040 29920 3052
rect 28767 3012 29920 3040
rect 28767 3009 28779 3012
rect 28721 3003 28779 3009
rect 29914 3000 29920 3012
rect 29972 3000 29978 3052
rect 30834 3040 30840 3052
rect 30024 3012 30840 3040
rect 25961 2975 26019 2981
rect 25961 2941 25973 2975
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 25976 2904 26004 2935
rect 26878 2932 26884 2984
rect 26936 2972 26942 2984
rect 28813 2975 28871 2981
rect 28813 2972 28825 2975
rect 26936 2944 28825 2972
rect 26936 2932 26942 2944
rect 28813 2941 28825 2944
rect 28859 2941 28871 2975
rect 30024 2972 30052 3012
rect 30834 3000 30840 3012
rect 30892 3000 30898 3052
rect 31113 3043 31171 3049
rect 31113 3009 31125 3043
rect 31159 3040 31171 3043
rect 31478 3040 31484 3052
rect 31159 3012 31484 3040
rect 31159 3009 31171 3012
rect 31113 3003 31171 3009
rect 31478 3000 31484 3012
rect 31536 3040 31542 3052
rect 34977 3043 35035 3049
rect 31536 3012 32996 3040
rect 31536 3000 31542 3012
rect 28813 2935 28871 2941
rect 28920 2944 30052 2972
rect 28920 2904 28948 2944
rect 30098 2932 30104 2984
rect 30156 2932 30162 2984
rect 30929 2975 30987 2981
rect 30929 2941 30941 2975
rect 30975 2972 30987 2975
rect 31662 2972 31668 2984
rect 30975 2944 31668 2972
rect 30975 2941 30987 2944
rect 30929 2935 30987 2941
rect 31662 2932 31668 2944
rect 31720 2932 31726 2984
rect 32214 2932 32220 2984
rect 32272 2932 32278 2984
rect 25976 2876 28948 2904
rect 29457 2907 29515 2913
rect 29457 2873 29469 2907
rect 29503 2904 29515 2907
rect 30006 2904 30012 2916
rect 29503 2876 30012 2904
rect 29503 2873 29515 2876
rect 29457 2867 29515 2873
rect 30006 2864 30012 2876
rect 30064 2864 30070 2916
rect 32968 2913 32996 3012
rect 34977 3009 34989 3043
rect 35023 3040 35035 3043
rect 35728 3040 35756 3080
rect 44910 3068 44916 3080
rect 44968 3068 44974 3120
rect 55140 3108 55168 3148
rect 57790 3136 57796 3148
rect 57848 3136 57854 3188
rect 57885 3179 57943 3185
rect 57885 3145 57897 3179
rect 57931 3176 57943 3179
rect 58986 3176 58992 3188
rect 57931 3148 58992 3176
rect 57931 3145 57943 3148
rect 57885 3139 57943 3145
rect 58986 3136 58992 3148
rect 59044 3136 59050 3188
rect 59078 3136 59084 3188
rect 59136 3136 59142 3188
rect 59541 3179 59599 3185
rect 59541 3145 59553 3179
rect 59587 3176 59599 3179
rect 62482 3176 62488 3188
rect 59587 3148 62488 3176
rect 59587 3145 59599 3148
rect 59541 3139 59599 3145
rect 62482 3136 62488 3148
rect 62540 3136 62546 3188
rect 63494 3136 63500 3188
rect 63552 3136 63558 3188
rect 66530 3136 66536 3188
rect 66588 3136 66594 3188
rect 69198 3136 69204 3188
rect 69256 3136 69262 3188
rect 59170 3108 59176 3120
rect 47780 3080 55168 3108
rect 55876 3080 59176 3108
rect 35023 3012 35756 3040
rect 35820 3012 37596 3040
rect 35023 3009 35035 3012
rect 34977 3003 35035 3009
rect 33134 2932 33140 2984
rect 33192 2972 33198 2984
rect 35820 2972 35848 3012
rect 33192 2944 35848 2972
rect 33192 2932 33198 2944
rect 35894 2932 35900 2984
rect 35952 2972 35958 2984
rect 36541 2975 36599 2981
rect 36541 2972 36553 2975
rect 35952 2944 36553 2972
rect 35952 2932 35958 2944
rect 36541 2941 36553 2944
rect 36587 2941 36599 2975
rect 36541 2935 36599 2941
rect 37458 2932 37464 2984
rect 37516 2932 37522 2984
rect 37568 2972 37596 3012
rect 37642 3000 37648 3052
rect 37700 3000 37706 3052
rect 38194 3040 38200 3052
rect 37752 3012 38200 3040
rect 37752 2972 37780 3012
rect 38194 3000 38200 3012
rect 38252 3000 38258 3052
rect 38378 3000 38384 3052
rect 38436 3000 38442 3052
rect 38838 3000 38844 3052
rect 38896 3000 38902 3052
rect 39114 3000 39120 3052
rect 39172 3000 39178 3052
rect 41322 3000 41328 3052
rect 41380 3000 41386 3052
rect 41601 3043 41659 3049
rect 41601 3009 41613 3043
rect 41647 3040 41659 3043
rect 41690 3040 41696 3052
rect 41647 3012 41696 3040
rect 41647 3009 41659 3012
rect 41601 3003 41659 3009
rect 41690 3000 41696 3012
rect 41748 3000 41754 3052
rect 42061 3043 42119 3049
rect 42061 3009 42073 3043
rect 42107 3040 42119 3043
rect 42426 3040 42432 3052
rect 42107 3012 42432 3040
rect 42107 3009 42119 3012
rect 42061 3003 42119 3009
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 43916 3012 44588 3040
rect 37568 2944 37780 2972
rect 37826 2932 37832 2984
rect 37884 2932 37890 2984
rect 37918 2932 37924 2984
rect 37976 2972 37982 2984
rect 40954 2972 40960 2984
rect 37976 2944 40960 2972
rect 37976 2932 37982 2944
rect 40954 2932 40960 2944
rect 41012 2932 41018 2984
rect 42242 2932 42248 2984
rect 42300 2972 42306 2984
rect 42337 2975 42395 2981
rect 42337 2972 42349 2975
rect 42300 2944 42349 2972
rect 42300 2932 42306 2944
rect 42337 2941 42349 2944
rect 42383 2941 42395 2975
rect 42337 2935 42395 2941
rect 32953 2907 33011 2913
rect 32953 2873 32965 2907
rect 32999 2904 33011 2907
rect 32999 2876 33548 2904
rect 32999 2873 33011 2876
rect 32953 2867 33011 2873
rect 27985 2839 28043 2845
rect 27985 2805 27997 2839
rect 28031 2836 28043 2839
rect 29086 2836 29092 2848
rect 28031 2808 29092 2836
rect 28031 2805 28043 2808
rect 27985 2799 28043 2805
rect 29086 2796 29092 2808
rect 29144 2796 29150 2848
rect 30285 2839 30343 2845
rect 30285 2805 30297 2839
rect 30331 2836 30343 2839
rect 30558 2836 30564 2848
rect 30331 2808 30564 2836
rect 30331 2805 30343 2808
rect 30285 2799 30343 2805
rect 30558 2796 30564 2808
rect 30616 2796 30622 2848
rect 31018 2796 31024 2848
rect 31076 2836 31082 2848
rect 31205 2839 31263 2845
rect 31205 2836 31217 2839
rect 31076 2808 31217 2836
rect 31076 2796 31082 2808
rect 31205 2805 31217 2808
rect 31251 2805 31263 2839
rect 31205 2799 31263 2805
rect 31294 2796 31300 2848
rect 31352 2836 31358 2848
rect 33134 2836 33140 2848
rect 31352 2808 33140 2836
rect 31352 2796 31358 2808
rect 33134 2796 33140 2808
rect 33192 2796 33198 2848
rect 33229 2839 33287 2845
rect 33229 2805 33241 2839
rect 33275 2836 33287 2839
rect 33410 2836 33416 2848
rect 33275 2808 33416 2836
rect 33275 2805 33287 2808
rect 33229 2799 33287 2805
rect 33410 2796 33416 2808
rect 33468 2796 33474 2848
rect 33520 2836 33548 2876
rect 35066 2864 35072 2916
rect 35124 2864 35130 2916
rect 43916 2904 43944 3012
rect 43993 2975 44051 2981
rect 43993 2941 44005 2975
rect 44039 2972 44051 2975
rect 44039 2944 44404 2972
rect 44039 2941 44051 2944
rect 43993 2935 44051 2941
rect 35176 2876 43944 2904
rect 35176 2836 35204 2876
rect 33520 2808 35204 2836
rect 35986 2796 35992 2848
rect 36044 2796 36050 2848
rect 36078 2796 36084 2848
rect 36136 2836 36142 2848
rect 42518 2836 42524 2848
rect 36136 2808 42524 2836
rect 36136 2796 36142 2808
rect 42518 2796 42524 2808
rect 42576 2796 42582 2848
rect 42978 2796 42984 2848
rect 43036 2796 43042 2848
rect 44376 2836 44404 2944
rect 44560 2904 44588 3012
rect 44634 3000 44640 3052
rect 44692 3000 44698 3052
rect 45002 3000 45008 3052
rect 45060 3040 45066 3052
rect 45177 3043 45235 3049
rect 45177 3040 45189 3043
rect 45060 3012 45189 3040
rect 45060 3000 45066 3012
rect 45177 3009 45189 3012
rect 45223 3009 45235 3043
rect 45177 3003 45235 3009
rect 46106 3000 46112 3052
rect 46164 3040 46170 3052
rect 47670 3040 47676 3052
rect 46164 3012 47676 3040
rect 46164 3000 46170 3012
rect 47670 3000 47676 3012
rect 47728 3000 47734 3052
rect 44913 2975 44971 2981
rect 44913 2941 44925 2975
rect 44959 2972 44971 2975
rect 47780 2972 47808 3080
rect 48038 3000 48044 3052
rect 48096 3040 48102 3052
rect 55876 3040 55904 3080
rect 59170 3068 59176 3080
rect 59228 3068 59234 3120
rect 60550 3068 60556 3120
rect 60608 3068 60614 3120
rect 62117 3111 62175 3117
rect 62117 3077 62129 3111
rect 62163 3108 62175 3111
rect 62298 3108 62304 3120
rect 62163 3080 62304 3108
rect 62163 3077 62175 3080
rect 62117 3071 62175 3077
rect 62298 3068 62304 3080
rect 62356 3068 62362 3120
rect 63586 3108 63592 3120
rect 62408 3080 63592 3108
rect 48096 3012 55904 3040
rect 58161 3043 58219 3049
rect 48096 3000 48102 3012
rect 58161 3009 58173 3043
rect 58207 3040 58219 3043
rect 59262 3040 59268 3052
rect 58207 3012 59268 3040
rect 58207 3009 58219 3012
rect 58161 3003 58219 3009
rect 59262 3000 59268 3012
rect 59320 3000 59326 3052
rect 59630 3000 59636 3052
rect 59688 3000 59694 3052
rect 61562 3000 61568 3052
rect 61620 3040 61626 3052
rect 62408 3040 62436 3080
rect 63586 3068 63592 3080
rect 63644 3068 63650 3120
rect 61620 3012 62436 3040
rect 61620 3000 61626 3012
rect 62666 3000 62672 3052
rect 62724 3040 62730 3052
rect 64601 3043 64659 3049
rect 64601 3040 64613 3043
rect 62724 3012 64613 3040
rect 62724 3000 62730 3012
rect 64601 3009 64613 3012
rect 64647 3009 64659 3043
rect 64601 3003 64659 3009
rect 69382 3000 69388 3052
rect 69440 3000 69446 3052
rect 44959 2944 47808 2972
rect 44959 2941 44971 2944
rect 44913 2935 44971 2941
rect 48130 2932 48136 2984
rect 48188 2972 48194 2984
rect 63862 2972 63868 2984
rect 48188 2944 63868 2972
rect 48188 2932 48194 2944
rect 63862 2932 63868 2944
rect 63920 2932 63926 2984
rect 63954 2932 63960 2984
rect 64012 2932 64018 2984
rect 64690 2932 64696 2984
rect 64748 2972 64754 2984
rect 65061 2975 65119 2981
rect 65061 2972 65073 2975
rect 64748 2944 65073 2972
rect 64748 2932 64754 2944
rect 65061 2941 65073 2944
rect 65107 2941 65119 2975
rect 65061 2935 65119 2941
rect 67177 2975 67235 2981
rect 67177 2941 67189 2975
rect 67223 2972 67235 2975
rect 67634 2972 67640 2984
rect 67223 2944 67640 2972
rect 67223 2941 67235 2944
rect 67177 2935 67235 2941
rect 67634 2932 67640 2944
rect 67692 2932 67698 2984
rect 68554 2932 68560 2984
rect 68612 2972 68618 2984
rect 69845 2975 69903 2981
rect 69845 2972 69857 2975
rect 68612 2944 69857 2972
rect 68612 2932 68618 2944
rect 69845 2941 69857 2944
rect 69891 2941 69903 2975
rect 69845 2935 69903 2941
rect 66438 2904 66444 2916
rect 44560 2876 66444 2904
rect 66438 2864 66444 2876
rect 66496 2864 66502 2916
rect 45094 2836 45100 2848
rect 44376 2808 45100 2836
rect 45094 2796 45100 2808
rect 45152 2796 45158 2848
rect 45462 2796 45468 2848
rect 45520 2836 45526 2848
rect 50798 2836 50804 2848
rect 45520 2808 50804 2836
rect 45520 2796 45526 2808
rect 50798 2796 50804 2808
rect 50856 2796 50862 2848
rect 59170 2796 59176 2848
rect 59228 2836 59234 2848
rect 62758 2836 62764 2848
rect 59228 2808 62764 2836
rect 59228 2796 59234 2808
rect 62758 2796 62764 2808
rect 62816 2796 62822 2848
rect 64509 2839 64567 2845
rect 64509 2805 64521 2839
rect 64555 2836 64567 2839
rect 65518 2836 65524 2848
rect 64555 2808 65524 2836
rect 64555 2805 64567 2808
rect 64509 2799 64567 2805
rect 65518 2796 65524 2808
rect 65576 2796 65582 2848
rect 67729 2839 67787 2845
rect 67729 2805 67741 2839
rect 67775 2836 67787 2839
rect 68094 2836 68100 2848
rect 67775 2808 68100 2836
rect 67775 2805 67787 2808
rect 67729 2799 67787 2805
rect 68094 2796 68100 2808
rect 68152 2796 68158 2848
rect 1012 2746 74980 2768
rect 1012 2694 1858 2746
rect 1910 2694 1922 2746
rect 1974 2694 1986 2746
rect 2038 2694 2050 2746
rect 2102 2694 2114 2746
rect 2166 2694 11858 2746
rect 11910 2694 11922 2746
rect 11974 2694 11986 2746
rect 12038 2694 12050 2746
rect 12102 2694 12114 2746
rect 12166 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 21986 2746
rect 22038 2694 22050 2746
rect 22102 2694 22114 2746
rect 22166 2694 31858 2746
rect 31910 2694 31922 2746
rect 31974 2694 31986 2746
rect 32038 2694 32050 2746
rect 32102 2694 32114 2746
rect 32166 2694 41858 2746
rect 41910 2694 41922 2746
rect 41974 2694 41986 2746
rect 42038 2694 42050 2746
rect 42102 2694 42114 2746
rect 42166 2694 51858 2746
rect 51910 2694 51922 2746
rect 51974 2694 51986 2746
rect 52038 2694 52050 2746
rect 52102 2694 52114 2746
rect 52166 2694 61858 2746
rect 61910 2694 61922 2746
rect 61974 2694 61986 2746
rect 62038 2694 62050 2746
rect 62102 2694 62114 2746
rect 62166 2694 71858 2746
rect 71910 2694 71922 2746
rect 71974 2694 71986 2746
rect 72038 2694 72050 2746
rect 72102 2694 72114 2746
rect 72166 2694 74980 2746
rect 1012 2672 74980 2694
rect 26697 2635 26755 2641
rect 26697 2601 26709 2635
rect 26743 2632 26755 2635
rect 27154 2632 27160 2644
rect 26743 2604 27160 2632
rect 26743 2601 26755 2604
rect 26697 2595 26755 2601
rect 27154 2592 27160 2604
rect 27212 2592 27218 2644
rect 29273 2635 29331 2641
rect 29273 2601 29285 2635
rect 29319 2632 29331 2635
rect 30098 2632 30104 2644
rect 29319 2604 30104 2632
rect 29319 2601 29331 2604
rect 29273 2595 29331 2601
rect 30098 2592 30104 2604
rect 30156 2592 30162 2644
rect 31389 2635 31447 2641
rect 31389 2601 31401 2635
rect 31435 2632 31447 2635
rect 32214 2632 32220 2644
rect 31435 2604 32220 2632
rect 31435 2601 31447 2604
rect 31389 2595 31447 2601
rect 32214 2592 32220 2604
rect 32272 2592 32278 2644
rect 33597 2635 33655 2641
rect 33597 2601 33609 2635
rect 33643 2632 33655 2635
rect 33870 2632 33876 2644
rect 33643 2604 33876 2632
rect 33643 2601 33655 2604
rect 33597 2595 33655 2601
rect 33870 2592 33876 2604
rect 33928 2592 33934 2644
rect 36354 2592 36360 2644
rect 36412 2632 36418 2644
rect 36633 2635 36691 2641
rect 36633 2632 36645 2635
rect 36412 2604 36645 2632
rect 36412 2592 36418 2604
rect 36633 2601 36645 2604
rect 36679 2601 36691 2635
rect 36633 2595 36691 2601
rect 37642 2592 37648 2644
rect 37700 2632 37706 2644
rect 37737 2635 37795 2641
rect 37737 2632 37749 2635
rect 37700 2604 37749 2632
rect 37700 2592 37706 2604
rect 37737 2601 37749 2604
rect 37783 2601 37795 2635
rect 37737 2595 37795 2601
rect 37826 2592 37832 2644
rect 37884 2592 37890 2644
rect 39114 2592 39120 2644
rect 39172 2632 39178 2644
rect 39393 2635 39451 2641
rect 39393 2632 39405 2635
rect 39172 2604 39405 2632
rect 39172 2592 39178 2604
rect 39393 2601 39405 2604
rect 39439 2601 39451 2635
rect 39393 2595 39451 2601
rect 41598 2592 41604 2644
rect 41656 2592 41662 2644
rect 41690 2592 41696 2644
rect 41748 2592 41754 2644
rect 42426 2592 42432 2644
rect 42484 2592 42490 2644
rect 44545 2635 44603 2641
rect 44545 2601 44557 2635
rect 44591 2632 44603 2635
rect 44634 2632 44640 2644
rect 44591 2604 44640 2632
rect 44591 2601 44603 2604
rect 44545 2595 44603 2601
rect 44634 2592 44640 2604
rect 44692 2592 44698 2644
rect 46017 2635 46075 2641
rect 46017 2601 46029 2635
rect 46063 2632 46075 2635
rect 52454 2632 52460 2644
rect 46063 2604 52460 2632
rect 46063 2601 46075 2604
rect 46017 2595 46075 2601
rect 52454 2592 52460 2604
rect 52512 2592 52518 2644
rect 52733 2635 52791 2641
rect 52733 2601 52745 2635
rect 52779 2632 52791 2635
rect 52779 2604 62804 2632
rect 52779 2601 52791 2604
rect 52733 2595 52791 2601
rect 29641 2567 29699 2573
rect 29641 2533 29653 2567
rect 29687 2564 29699 2567
rect 48406 2564 48412 2576
rect 29687 2536 48412 2564
rect 29687 2533 29699 2536
rect 29641 2527 29699 2533
rect 48406 2524 48412 2536
rect 48464 2524 48470 2576
rect 48685 2567 48743 2573
rect 48685 2533 48697 2567
rect 48731 2533 48743 2567
rect 48685 2527 48743 2533
rect 25961 2499 26019 2505
rect 25961 2465 25973 2499
rect 26007 2496 26019 2499
rect 26234 2496 26240 2508
rect 26007 2468 26240 2496
rect 26007 2465 26019 2468
rect 25961 2459 26019 2465
rect 26234 2456 26240 2468
rect 26292 2456 26298 2508
rect 27062 2456 27068 2508
rect 27120 2496 27126 2508
rect 27120 2468 28994 2496
rect 27120 2456 27126 2468
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 24949 2431 25007 2437
rect 24949 2428 24961 2431
rect 24912 2400 24961 2428
rect 24912 2388 24918 2400
rect 24949 2397 24961 2400
rect 24995 2397 25007 2431
rect 24949 2391 25007 2397
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2428 26203 2431
rect 27154 2428 27160 2440
rect 26191 2400 27160 2428
rect 26191 2397 26203 2400
rect 26145 2391 26203 2397
rect 27154 2388 27160 2400
rect 27212 2388 27218 2440
rect 28166 2388 28172 2440
rect 28224 2388 28230 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2397 28411 2431
rect 28353 2391 28411 2397
rect 28721 2431 28779 2437
rect 28721 2397 28733 2431
rect 28767 2397 28779 2431
rect 28966 2428 28994 2468
rect 30558 2456 30564 2508
rect 30616 2456 30622 2508
rect 32490 2496 32496 2508
rect 30668 2468 32496 2496
rect 30668 2428 30696 2468
rect 32490 2456 32496 2468
rect 32548 2456 32554 2508
rect 33594 2456 33600 2508
rect 33652 2496 33658 2508
rect 34241 2499 34299 2505
rect 34241 2496 34253 2499
rect 33652 2468 34253 2496
rect 33652 2456 33658 2468
rect 34241 2465 34253 2468
rect 34287 2465 34299 2499
rect 34241 2459 34299 2465
rect 34348 2468 35756 2496
rect 28966 2400 30696 2428
rect 28721 2391 28779 2397
rect 26786 2320 26792 2372
rect 26844 2360 26850 2372
rect 26973 2363 27031 2369
rect 26973 2360 26985 2363
rect 26844 2332 26985 2360
rect 26844 2320 26850 2332
rect 26973 2329 26985 2332
rect 27019 2329 27031 2363
rect 26973 2323 27031 2329
rect 27614 2320 27620 2372
rect 27672 2360 27678 2372
rect 28368 2360 28396 2391
rect 27672 2332 28396 2360
rect 27672 2320 27678 2332
rect 25130 2252 25136 2304
rect 25188 2252 25194 2304
rect 25222 2252 25228 2304
rect 25280 2292 25286 2304
rect 25317 2295 25375 2301
rect 25317 2292 25329 2295
rect 25280 2264 25329 2292
rect 25280 2252 25286 2264
rect 25317 2261 25329 2264
rect 25363 2261 25375 2295
rect 25317 2255 25375 2261
rect 28442 2252 28448 2304
rect 28500 2252 28506 2304
rect 28736 2292 28764 2391
rect 30834 2388 30840 2440
rect 30892 2388 30898 2440
rect 31478 2388 31484 2440
rect 31536 2388 31542 2440
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33045 2431 33103 2437
rect 33045 2397 33057 2431
rect 33091 2428 33103 2431
rect 33689 2431 33747 2437
rect 33689 2428 33701 2431
rect 33091 2400 33701 2428
rect 33091 2397 33103 2400
rect 33045 2391 33103 2397
rect 33689 2397 33701 2400
rect 33735 2397 33747 2431
rect 33689 2391 33747 2397
rect 29825 2363 29883 2369
rect 29825 2329 29837 2363
rect 29871 2360 29883 2363
rect 30009 2363 30067 2369
rect 30009 2360 30021 2363
rect 29871 2332 30021 2360
rect 29871 2329 29883 2332
rect 29825 2323 29883 2329
rect 30009 2329 30021 2332
rect 30055 2329 30067 2363
rect 32324 2360 32352 2391
rect 33962 2388 33968 2440
rect 34020 2428 34026 2440
rect 34348 2428 34376 2468
rect 34020 2400 34376 2428
rect 34020 2388 34026 2400
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35621 2431 35679 2437
rect 35621 2428 35633 2431
rect 35032 2400 35633 2428
rect 35032 2388 35038 2400
rect 35621 2397 35633 2400
rect 35667 2397 35679 2431
rect 35621 2391 35679 2397
rect 35069 2363 35127 2369
rect 35069 2360 35081 2363
rect 32324 2332 35081 2360
rect 30009 2323 30067 2329
rect 35069 2329 35081 2332
rect 35115 2329 35127 2363
rect 35069 2323 35127 2329
rect 31294 2292 31300 2304
rect 28736 2264 31300 2292
rect 31294 2252 31300 2264
rect 31352 2252 31358 2304
rect 32125 2295 32183 2301
rect 32125 2261 32137 2295
rect 32171 2292 32183 2295
rect 32490 2292 32496 2304
rect 32171 2264 32496 2292
rect 32171 2261 32183 2264
rect 32125 2255 32183 2261
rect 32490 2252 32496 2264
rect 32548 2252 32554 2304
rect 32861 2295 32919 2301
rect 32861 2261 32873 2295
rect 32907 2292 32919 2295
rect 35158 2292 35164 2304
rect 32907 2264 35164 2292
rect 32907 2261 32919 2264
rect 32861 2255 32919 2261
rect 35158 2252 35164 2264
rect 35216 2252 35222 2304
rect 35728 2292 35756 2468
rect 35986 2456 35992 2508
rect 36044 2456 36050 2508
rect 42978 2456 42984 2508
rect 43036 2456 43042 2508
rect 48700 2496 48728 2527
rect 51626 2524 51632 2576
rect 51684 2564 51690 2576
rect 57333 2567 57391 2573
rect 51684 2536 57192 2564
rect 51684 2524 51690 2536
rect 56686 2496 56692 2508
rect 48700 2468 51028 2496
rect 36998 2388 37004 2440
rect 37056 2428 37062 2440
rect 37093 2431 37151 2437
rect 37093 2428 37105 2431
rect 37056 2400 37105 2428
rect 37056 2388 37062 2400
rect 37093 2397 37105 2400
rect 37139 2397 37151 2431
rect 37093 2391 37151 2397
rect 37734 2388 37740 2440
rect 37792 2428 37798 2440
rect 38381 2431 38439 2437
rect 38381 2428 38393 2431
rect 37792 2400 38393 2428
rect 37792 2388 37798 2400
rect 38381 2397 38393 2400
rect 38427 2397 38439 2431
rect 38381 2391 38439 2397
rect 38746 2388 38752 2440
rect 38804 2388 38810 2440
rect 40589 2431 40647 2437
rect 40589 2397 40601 2431
rect 40635 2428 40647 2431
rect 40678 2428 40684 2440
rect 40635 2400 40684 2428
rect 40635 2397 40647 2400
rect 40589 2391 40647 2397
rect 40678 2388 40684 2400
rect 40736 2388 40742 2440
rect 41049 2431 41107 2437
rect 41049 2397 41061 2431
rect 41095 2428 41107 2431
rect 41414 2428 41420 2440
rect 41095 2400 41420 2428
rect 41095 2397 41107 2400
rect 41049 2391 41107 2397
rect 41414 2388 41420 2400
rect 41472 2388 41478 2440
rect 42337 2431 42395 2437
rect 42337 2397 42349 2431
rect 42383 2428 42395 2431
rect 42702 2428 42708 2440
rect 42383 2400 42708 2428
rect 42383 2397 42395 2400
rect 42337 2391 42395 2397
rect 42702 2388 42708 2400
rect 42760 2388 42766 2440
rect 42794 2388 42800 2440
rect 42852 2428 42858 2440
rect 43165 2431 43223 2437
rect 43165 2428 43177 2431
rect 42852 2400 43177 2428
rect 42852 2388 42858 2400
rect 43165 2397 43177 2400
rect 43211 2397 43223 2431
rect 43165 2391 43223 2397
rect 43809 2431 43867 2437
rect 43809 2397 43821 2431
rect 43855 2428 43867 2431
rect 43901 2431 43959 2437
rect 43901 2428 43913 2431
rect 43855 2400 43913 2428
rect 43855 2397 43867 2400
rect 43809 2391 43867 2397
rect 43901 2397 43913 2400
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 45189 2431 45247 2437
rect 45189 2397 45201 2431
rect 45235 2428 45247 2431
rect 45462 2428 45468 2440
rect 45235 2400 45468 2428
rect 45235 2397 45247 2400
rect 45189 2391 45247 2397
rect 45462 2388 45468 2400
rect 45520 2388 45526 2440
rect 45741 2431 45799 2437
rect 45741 2397 45753 2431
rect 45787 2428 45799 2431
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 45787 2400 45845 2428
rect 45787 2397 45799 2400
rect 45741 2391 45799 2397
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 46477 2431 46535 2437
rect 46477 2397 46489 2431
rect 46523 2428 46535 2431
rect 46934 2428 46940 2440
rect 46523 2400 46940 2428
rect 46523 2397 46535 2400
rect 46477 2391 46535 2397
rect 46934 2388 46940 2400
rect 46992 2388 46998 2440
rect 47394 2388 47400 2440
rect 47452 2428 47458 2440
rect 47489 2431 47547 2437
rect 47489 2428 47501 2431
rect 47452 2400 47501 2428
rect 47452 2388 47458 2400
rect 47489 2397 47501 2400
rect 47535 2397 47547 2431
rect 47489 2391 47547 2397
rect 48869 2431 48927 2437
rect 48869 2397 48881 2431
rect 48915 2428 48927 2431
rect 48961 2431 49019 2437
rect 48961 2428 48973 2431
rect 48915 2400 48973 2428
rect 48915 2397 48927 2400
rect 48869 2391 48927 2397
rect 48961 2397 48973 2400
rect 49007 2397 49019 2431
rect 48961 2391 49019 2397
rect 49418 2388 49424 2440
rect 49476 2428 49482 2440
rect 49513 2431 49571 2437
rect 49513 2428 49525 2431
rect 49476 2400 49525 2428
rect 49476 2388 49482 2400
rect 49513 2397 49525 2400
rect 49559 2397 49571 2431
rect 49513 2391 49571 2397
rect 50154 2388 50160 2440
rect 50212 2388 50218 2440
rect 51000 2428 51028 2468
rect 51644 2468 56692 2496
rect 51644 2428 51672 2468
rect 56686 2456 56692 2468
rect 56744 2456 56750 2508
rect 51000 2400 51672 2428
rect 51721 2431 51779 2437
rect 51721 2397 51733 2431
rect 51767 2428 51779 2431
rect 52638 2428 52644 2440
rect 51767 2400 52644 2428
rect 51767 2397 51779 2400
rect 51721 2391 51779 2397
rect 52638 2388 52644 2400
rect 52696 2388 52702 2440
rect 53650 2388 53656 2440
rect 53708 2388 53714 2440
rect 55309 2431 55367 2437
rect 55309 2397 55321 2431
rect 55355 2428 55367 2431
rect 55582 2428 55588 2440
rect 55355 2400 55588 2428
rect 55355 2397 55367 2400
rect 55309 2391 55367 2397
rect 55582 2388 55588 2400
rect 55640 2388 55646 2440
rect 56318 2388 56324 2440
rect 56376 2388 56382 2440
rect 40313 2363 40371 2369
rect 40313 2329 40325 2363
rect 40359 2360 40371 2363
rect 51626 2360 51632 2372
rect 40359 2332 51632 2360
rect 40359 2329 40371 2332
rect 40313 2323 40371 2329
rect 51626 2320 51632 2332
rect 51684 2320 51690 2372
rect 52273 2363 52331 2369
rect 52273 2329 52285 2363
rect 52319 2360 52331 2363
rect 52457 2363 52515 2369
rect 52457 2360 52469 2363
rect 52319 2332 52469 2360
rect 52319 2329 52331 2332
rect 52273 2323 52331 2329
rect 52457 2329 52469 2332
rect 52503 2329 52515 2363
rect 52457 2323 52515 2329
rect 54205 2363 54263 2369
rect 54205 2329 54217 2363
rect 54251 2360 54263 2363
rect 54389 2363 54447 2369
rect 54389 2360 54401 2363
rect 54251 2332 54401 2360
rect 54251 2329 54263 2332
rect 54205 2323 54263 2329
rect 54389 2329 54401 2332
rect 54435 2329 54447 2363
rect 54389 2323 54447 2329
rect 54757 2363 54815 2369
rect 54757 2329 54769 2363
rect 54803 2360 54815 2363
rect 56873 2363 56931 2369
rect 54803 2332 56824 2360
rect 54803 2329 54815 2332
rect 54757 2323 54815 2329
rect 46842 2292 46848 2304
rect 35728 2264 46848 2292
rect 46842 2252 46848 2264
rect 46900 2252 46906 2304
rect 47026 2252 47032 2304
rect 47084 2252 47090 2304
rect 48130 2252 48136 2304
rect 48188 2252 48194 2304
rect 50798 2252 50804 2304
rect 50856 2252 50862 2304
rect 55766 2252 55772 2304
rect 55824 2292 55830 2304
rect 55861 2295 55919 2301
rect 55861 2292 55873 2295
rect 55824 2264 55873 2292
rect 55824 2252 55830 2264
rect 55861 2261 55873 2264
rect 55907 2261 55919 2295
rect 56796 2292 56824 2332
rect 56873 2329 56885 2363
rect 56919 2360 56931 2363
rect 57057 2363 57115 2369
rect 57057 2360 57069 2363
rect 56919 2332 57069 2360
rect 56919 2329 56931 2332
rect 56873 2323 56931 2329
rect 57057 2329 57069 2332
rect 57103 2329 57115 2363
rect 57164 2360 57192 2536
rect 57333 2533 57345 2567
rect 57379 2564 57391 2567
rect 62666 2564 62672 2576
rect 57379 2536 62672 2564
rect 57379 2533 57391 2536
rect 57333 2527 57391 2533
rect 62666 2524 62672 2536
rect 62724 2524 62730 2576
rect 62776 2564 62804 2604
rect 63494 2592 63500 2644
rect 63552 2592 63558 2644
rect 65886 2592 65892 2644
rect 65944 2632 65950 2644
rect 66165 2635 66223 2641
rect 66165 2632 66177 2635
rect 65944 2604 66177 2632
rect 65944 2592 65950 2604
rect 66165 2601 66177 2604
rect 66211 2601 66223 2635
rect 66165 2595 66223 2601
rect 66530 2592 66536 2644
rect 66588 2592 66594 2644
rect 69198 2592 69204 2644
rect 69256 2592 69262 2644
rect 63770 2564 63776 2576
rect 62776 2536 63776 2564
rect 63770 2524 63776 2536
rect 63828 2524 63834 2576
rect 57514 2456 57520 2508
rect 57572 2496 57578 2508
rect 58069 2499 58127 2505
rect 58069 2496 58081 2499
rect 57572 2468 58081 2496
rect 57572 2456 57578 2468
rect 58069 2465 58081 2468
rect 58115 2465 58127 2499
rect 58069 2459 58127 2465
rect 59078 2456 59084 2508
rect 59136 2456 59142 2508
rect 60550 2456 60556 2508
rect 60608 2456 60614 2508
rect 61654 2456 61660 2508
rect 61712 2496 61718 2508
rect 64141 2499 64199 2505
rect 61712 2468 63724 2496
rect 61712 2456 61718 2468
rect 57422 2388 57428 2440
rect 57480 2428 57486 2440
rect 57609 2431 57667 2437
rect 57609 2428 57621 2431
rect 57480 2400 57621 2428
rect 57480 2388 57486 2400
rect 57609 2397 57621 2400
rect 57655 2397 57667 2431
rect 57609 2391 57667 2397
rect 58526 2388 58532 2440
rect 58584 2428 58590 2440
rect 59265 2431 59323 2437
rect 59265 2428 59277 2431
rect 58584 2400 59277 2428
rect 58584 2388 58590 2400
rect 59265 2397 59277 2400
rect 59311 2397 59323 2431
rect 59265 2391 59323 2397
rect 61378 2388 61384 2440
rect 61436 2428 61442 2440
rect 61841 2431 61899 2437
rect 61841 2428 61853 2431
rect 61436 2400 61853 2428
rect 61436 2388 61442 2400
rect 61841 2397 61853 2400
rect 61887 2397 61899 2431
rect 61841 2391 61899 2397
rect 62298 2388 62304 2440
rect 62356 2388 62362 2440
rect 63696 2437 63724 2468
rect 64141 2465 64153 2499
rect 64187 2465 64199 2499
rect 64141 2459 64199 2465
rect 63681 2431 63739 2437
rect 63681 2397 63693 2431
rect 63727 2397 63739 2431
rect 63681 2391 63739 2397
rect 60090 2360 60096 2372
rect 57164 2332 60096 2360
rect 57057 2323 57115 2329
rect 60090 2320 60096 2332
rect 60148 2320 60154 2372
rect 61105 2363 61163 2369
rect 61105 2329 61117 2363
rect 61151 2360 61163 2363
rect 61289 2363 61347 2369
rect 61289 2360 61301 2363
rect 61151 2332 61301 2360
rect 61151 2329 61163 2332
rect 61105 2323 61163 2329
rect 61289 2329 61301 2332
rect 61335 2329 61347 2363
rect 64156 2360 64184 2459
rect 65518 2456 65524 2508
rect 65576 2456 65582 2508
rect 65794 2456 65800 2508
rect 65852 2496 65858 2508
rect 67085 2499 67143 2505
rect 67085 2496 67097 2499
rect 65852 2468 67097 2496
rect 65852 2456 65858 2468
rect 67085 2465 67097 2468
rect 67131 2465 67143 2499
rect 67085 2459 67143 2465
rect 68370 2456 68376 2508
rect 68428 2456 68434 2508
rect 69842 2456 69848 2508
rect 69900 2496 69906 2508
rect 71593 2499 71651 2505
rect 71593 2496 71605 2499
rect 69900 2468 71605 2496
rect 69900 2456 69906 2468
rect 71593 2465 71605 2468
rect 71639 2465 71651 2499
rect 71593 2459 71651 2465
rect 65334 2388 65340 2440
rect 65392 2428 65398 2440
rect 66625 2431 66683 2437
rect 66625 2428 66637 2431
rect 65392 2400 66637 2428
rect 65392 2388 65398 2400
rect 66625 2397 66637 2400
rect 66671 2397 66683 2431
rect 66625 2391 66683 2397
rect 68094 2388 68100 2440
rect 68152 2388 68158 2440
rect 69474 2388 69480 2440
rect 69532 2388 69538 2440
rect 70670 2388 70676 2440
rect 70728 2388 70734 2440
rect 71317 2431 71375 2437
rect 71317 2397 71329 2431
rect 71363 2428 71375 2431
rect 71409 2431 71467 2437
rect 71409 2428 71421 2431
rect 71363 2400 71421 2428
rect 71363 2397 71375 2400
rect 71317 2391 71375 2397
rect 71409 2397 71421 2400
rect 71455 2397 71467 2431
rect 71409 2391 71467 2397
rect 72602 2388 72608 2440
rect 72660 2388 72666 2440
rect 61289 2323 61347 2329
rect 62040 2332 64184 2360
rect 59170 2292 59176 2304
rect 56796 2264 59176 2292
rect 55861 2255 55919 2261
rect 59170 2252 59176 2264
rect 59228 2252 59234 2304
rect 59909 2295 59967 2301
rect 59909 2261 59921 2295
rect 59955 2292 59967 2295
rect 59998 2292 60004 2304
rect 59955 2264 60004 2292
rect 59955 2261 59967 2264
rect 59909 2255 59967 2261
rect 59998 2252 60004 2264
rect 60056 2252 60062 2304
rect 61010 2252 61016 2304
rect 61068 2252 61074 2304
rect 61654 2252 61660 2304
rect 61712 2292 61718 2304
rect 62040 2292 62068 2332
rect 69658 2320 69664 2372
rect 69716 2360 69722 2372
rect 72329 2363 72387 2369
rect 72329 2360 72341 2363
rect 69716 2332 72341 2360
rect 69716 2320 69722 2332
rect 72329 2329 72341 2332
rect 72375 2329 72387 2363
rect 72329 2323 72387 2329
rect 61712 2264 62068 2292
rect 62117 2295 62175 2301
rect 61712 2252 61718 2264
rect 62117 2261 62129 2295
rect 62163 2292 62175 2295
rect 62390 2292 62396 2304
rect 62163 2264 62396 2292
rect 62163 2261 62175 2264
rect 62117 2255 62175 2261
rect 62390 2252 62396 2264
rect 62448 2252 62454 2304
rect 62574 2252 62580 2304
rect 62632 2292 62638 2304
rect 62853 2295 62911 2301
rect 62853 2292 62865 2295
rect 62632 2264 62865 2292
rect 62632 2252 62638 2264
rect 62853 2261 62865 2264
rect 62899 2261 62911 2295
rect 62853 2255 62911 2261
rect 63126 2252 63132 2304
rect 63184 2292 63190 2304
rect 64598 2292 64604 2304
rect 63184 2264 64604 2292
rect 63184 2252 63190 2264
rect 64598 2252 64604 2264
rect 64656 2252 64662 2304
rect 70029 2295 70087 2301
rect 70029 2261 70041 2295
rect 70075 2292 70087 2295
rect 70854 2292 70860 2304
rect 70075 2264 70860 2292
rect 70075 2261 70087 2264
rect 70029 2255 70087 2261
rect 70854 2252 70860 2264
rect 70912 2252 70918 2304
rect 1012 2202 74980 2224
rect 1012 2150 4210 2202
rect 4262 2150 4274 2202
rect 4326 2150 4338 2202
rect 4390 2150 4402 2202
rect 4454 2150 4466 2202
rect 4518 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 24466 2202
rect 24518 2150 34210 2202
rect 34262 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 44210 2202
rect 44262 2150 44274 2202
rect 44326 2150 44338 2202
rect 44390 2150 44402 2202
rect 44454 2150 44466 2202
rect 44518 2150 54210 2202
rect 54262 2150 54274 2202
rect 54326 2150 54338 2202
rect 54390 2150 54402 2202
rect 54454 2150 54466 2202
rect 54518 2150 64210 2202
rect 64262 2150 64274 2202
rect 64326 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 74210 2202
rect 74262 2150 74274 2202
rect 74326 2150 74338 2202
rect 74390 2150 74402 2202
rect 74454 2150 74466 2202
rect 74518 2150 74980 2202
rect 1012 2128 74980 2150
rect 24397 2091 24455 2097
rect 24397 2057 24409 2091
rect 24443 2057 24455 2091
rect 24397 2051 24455 2057
rect 25225 2091 25283 2097
rect 25225 2057 25237 2091
rect 25271 2088 25283 2091
rect 25682 2088 25688 2100
rect 25271 2060 25688 2088
rect 25271 2057 25283 2060
rect 25225 2051 25283 2057
rect 24412 2020 24440 2051
rect 25682 2048 25688 2060
rect 25740 2048 25746 2100
rect 25961 2091 26019 2097
rect 25961 2057 25973 2091
rect 26007 2088 26019 2091
rect 26602 2088 26608 2100
rect 26007 2060 26608 2088
rect 26007 2057 26019 2060
rect 25961 2051 26019 2057
rect 26602 2048 26608 2060
rect 26660 2048 26666 2100
rect 26694 2048 26700 2100
rect 26752 2048 26758 2100
rect 27062 2048 27068 2100
rect 27120 2048 27126 2100
rect 28442 2048 28448 2100
rect 28500 2088 28506 2100
rect 34054 2088 34060 2100
rect 28500 2060 34060 2088
rect 28500 2048 28506 2060
rect 34054 2048 34060 2060
rect 34112 2048 34118 2100
rect 36265 2091 36323 2097
rect 36265 2057 36277 2091
rect 36311 2088 36323 2091
rect 36538 2088 36544 2100
rect 36311 2060 36544 2088
rect 36311 2057 36323 2060
rect 36265 2051 36323 2057
rect 36538 2048 36544 2060
rect 36596 2048 36602 2100
rect 36998 2048 37004 2100
rect 37056 2048 37062 2100
rect 40678 2048 40684 2100
rect 40736 2048 40742 2100
rect 41414 2048 41420 2100
rect 41472 2048 41478 2100
rect 41690 2048 41696 2100
rect 41748 2088 41754 2100
rect 44726 2088 44732 2100
rect 41748 2060 44732 2088
rect 41748 2048 41754 2060
rect 44726 2048 44732 2060
rect 44784 2048 44790 2100
rect 45094 2048 45100 2100
rect 45152 2088 45158 2100
rect 45373 2091 45431 2097
rect 45373 2088 45385 2091
rect 45152 2060 45385 2088
rect 45152 2048 45158 2060
rect 45373 2057 45385 2060
rect 45419 2057 45431 2091
rect 45373 2051 45431 2057
rect 46934 2048 46940 2100
rect 46992 2048 46998 2100
rect 47578 2048 47584 2100
rect 47636 2048 47642 2100
rect 49418 2048 49424 2100
rect 49476 2048 49482 2100
rect 50433 2091 50491 2097
rect 50433 2057 50445 2091
rect 50479 2088 50491 2091
rect 50479 2060 51074 2088
rect 50479 2057 50491 2060
rect 50433 2051 50491 2057
rect 30193 2023 30251 2029
rect 24412 1992 30144 2020
rect 24213 1955 24271 1961
rect 24213 1921 24225 1955
rect 24259 1952 24271 1955
rect 24670 1952 24676 1964
rect 24259 1924 24676 1952
rect 24259 1921 24271 1924
rect 24213 1915 24271 1921
rect 24670 1912 24676 1924
rect 24728 1912 24734 1964
rect 25314 1912 25320 1964
rect 25372 1952 25378 1964
rect 26881 1955 26939 1961
rect 26881 1952 26893 1955
rect 25372 1924 26893 1952
rect 25372 1912 25378 1924
rect 26881 1921 26893 1924
rect 26927 1921 26939 1955
rect 26881 1915 26939 1921
rect 27433 1955 27491 1961
rect 27433 1921 27445 1955
rect 27479 1952 27491 1955
rect 27798 1952 27804 1964
rect 27479 1924 27804 1952
rect 27479 1921 27491 1924
rect 27433 1915 27491 1921
rect 27798 1912 27804 1924
rect 27856 1912 27862 1964
rect 29086 1912 29092 1964
rect 29144 1912 29150 1964
rect 30116 1952 30144 1992
rect 30193 1989 30205 2023
rect 30239 2020 30251 2023
rect 33962 2020 33968 2032
rect 30239 1992 33968 2020
rect 30239 1989 30251 1992
rect 30193 1983 30251 1989
rect 33962 1980 33968 1992
rect 34020 1980 34026 2032
rect 34882 1980 34888 2032
rect 34940 2020 34946 2032
rect 41138 2020 41144 2032
rect 34940 1992 41144 2020
rect 34940 1980 34946 1992
rect 41138 1980 41144 1992
rect 41196 1980 41202 2032
rect 48774 1980 48780 2032
rect 48832 2020 48838 2032
rect 51046 2020 51074 2060
rect 52638 2048 52644 2100
rect 52696 2048 52702 2100
rect 55582 2048 55588 2100
rect 55640 2048 55646 2100
rect 59078 2048 59084 2100
rect 59136 2048 59142 2100
rect 59449 2091 59507 2097
rect 59449 2057 59461 2091
rect 59495 2088 59507 2091
rect 59630 2088 59636 2100
rect 59495 2060 59636 2088
rect 59495 2057 59507 2060
rect 59449 2051 59507 2057
rect 59630 2048 59636 2060
rect 59688 2048 59694 2100
rect 60550 2048 60556 2100
rect 60608 2048 60614 2100
rect 61378 2048 61384 2100
rect 61436 2048 61442 2100
rect 66346 2088 66352 2100
rect 61488 2060 66352 2088
rect 61488 2020 61516 2060
rect 66346 2048 66352 2060
rect 66404 2048 66410 2100
rect 66530 2048 66536 2100
rect 66588 2048 66594 2100
rect 66990 2048 66996 2100
rect 67048 2088 67054 2100
rect 69109 2091 69167 2097
rect 67048 2060 68784 2088
rect 67048 2048 67054 2060
rect 48832 1992 50752 2020
rect 51046 1992 61516 2020
rect 62117 2023 62175 2029
rect 48832 1980 48838 1992
rect 31110 1952 31116 1964
rect 30116 1924 31116 1952
rect 31110 1912 31116 1924
rect 31168 1912 31174 1964
rect 31849 1955 31907 1961
rect 31849 1921 31861 1955
rect 31895 1952 31907 1955
rect 33042 1952 33048 1964
rect 31895 1924 33048 1952
rect 31895 1921 31907 1924
rect 31849 1915 31907 1921
rect 33042 1912 33048 1924
rect 33100 1912 33106 1964
rect 33502 1912 33508 1964
rect 33560 1912 33566 1964
rect 33870 1912 33876 1964
rect 33928 1952 33934 1964
rect 34149 1955 34207 1961
rect 34149 1952 34161 1955
rect 33928 1924 34161 1952
rect 33928 1912 33934 1924
rect 34149 1921 34161 1924
rect 34195 1921 34207 1955
rect 34149 1915 34207 1921
rect 34606 1912 34612 1964
rect 34664 1952 34670 1964
rect 37185 1955 37243 1961
rect 37185 1952 37197 1955
rect 34664 1924 37197 1952
rect 34664 1912 34670 1924
rect 37185 1921 37197 1924
rect 37231 1921 37243 1955
rect 37185 1915 37243 1921
rect 39025 1955 39083 1961
rect 39025 1921 39037 1955
rect 39071 1952 39083 1955
rect 39209 1955 39267 1961
rect 39209 1952 39221 1955
rect 39071 1924 39221 1952
rect 39071 1921 39083 1924
rect 39025 1915 39083 1921
rect 39209 1921 39221 1924
rect 39255 1921 39267 1955
rect 40497 1955 40555 1961
rect 40497 1952 40509 1955
rect 39209 1915 39267 1921
rect 39316 1924 40509 1952
rect 24581 1887 24639 1893
rect 24581 1853 24593 1887
rect 24627 1884 24639 1887
rect 25222 1884 25228 1896
rect 24627 1856 25228 1884
rect 24627 1853 24639 1856
rect 24581 1847 24639 1853
rect 25222 1844 25228 1856
rect 25280 1844 25286 1896
rect 25406 1844 25412 1896
rect 25464 1844 25470 1896
rect 26145 1887 26203 1893
rect 26145 1853 26157 1887
rect 26191 1884 26203 1887
rect 27522 1884 27528 1896
rect 26191 1856 27528 1884
rect 26191 1853 26203 1856
rect 26145 1847 26203 1853
rect 27522 1844 27528 1856
rect 27580 1844 27586 1896
rect 28445 1887 28503 1893
rect 28445 1853 28457 1887
rect 28491 1853 28503 1887
rect 28445 1847 28503 1853
rect 28460 1816 28488 1847
rect 30374 1844 30380 1896
rect 30432 1884 30438 1896
rect 30653 1887 30711 1893
rect 30653 1884 30665 1887
rect 30432 1856 30665 1884
rect 30432 1844 30438 1856
rect 30653 1853 30665 1856
rect 30699 1853 30711 1887
rect 30653 1847 30711 1853
rect 32214 1844 32220 1896
rect 32272 1884 32278 1896
rect 32493 1887 32551 1893
rect 32493 1884 32505 1887
rect 32272 1856 32505 1884
rect 32272 1844 32278 1856
rect 32493 1853 32505 1856
rect 32539 1853 32551 1887
rect 32493 1847 32551 1853
rect 34054 1844 34060 1896
rect 34112 1884 34118 1896
rect 34701 1887 34759 1893
rect 34701 1884 34713 1887
rect 34112 1856 34713 1884
rect 34112 1844 34118 1856
rect 34701 1853 34713 1856
rect 34747 1853 34759 1887
rect 34701 1847 34759 1853
rect 35618 1844 35624 1896
rect 35676 1844 35682 1896
rect 36449 1887 36507 1893
rect 36449 1853 36461 1887
rect 36495 1884 36507 1887
rect 37274 1884 37280 1896
rect 36495 1856 37280 1884
rect 36495 1853 36507 1856
rect 36449 1847 36507 1853
rect 37274 1844 37280 1856
rect 37332 1844 37338 1896
rect 37645 1887 37703 1893
rect 37645 1853 37657 1887
rect 37691 1853 37703 1887
rect 37645 1847 37703 1853
rect 28460 1788 36584 1816
rect 28166 1708 28172 1760
rect 28224 1748 28230 1760
rect 30558 1748 30564 1760
rect 28224 1720 30564 1748
rect 28224 1708 28230 1720
rect 30558 1708 30564 1720
rect 30616 1708 30622 1760
rect 32490 1708 32496 1760
rect 32548 1748 32554 1760
rect 35802 1748 35808 1760
rect 32548 1720 35808 1748
rect 32548 1708 32554 1720
rect 35802 1708 35808 1720
rect 35860 1708 35866 1760
rect 36556 1748 36584 1788
rect 36814 1776 36820 1828
rect 36872 1816 36878 1828
rect 37660 1816 37688 1847
rect 39114 1844 39120 1896
rect 39172 1884 39178 1896
rect 39316 1884 39344 1924
rect 40497 1921 40509 1924
rect 40543 1921 40555 1955
rect 40497 1915 40555 1921
rect 41230 1912 41236 1964
rect 41288 1912 41294 1964
rect 41414 1912 41420 1964
rect 41472 1952 41478 1964
rect 41969 1955 42027 1961
rect 41969 1952 41981 1955
rect 41472 1924 41981 1952
rect 41472 1912 41478 1924
rect 41969 1921 41981 1924
rect 42015 1921 42027 1955
rect 41969 1915 42027 1921
rect 42429 1955 42487 1961
rect 42429 1921 42441 1955
rect 42475 1921 42487 1955
rect 42429 1915 42487 1921
rect 39172 1856 39344 1884
rect 39853 1887 39911 1893
rect 39172 1844 39178 1856
rect 39853 1853 39865 1887
rect 39899 1884 39911 1887
rect 39945 1887 40003 1893
rect 39945 1884 39957 1887
rect 39899 1856 39957 1884
rect 39899 1853 39911 1856
rect 39853 1847 39911 1853
rect 39945 1853 39957 1856
rect 39991 1853 40003 1887
rect 39945 1847 40003 1853
rect 40034 1844 40040 1896
rect 40092 1884 40098 1896
rect 42444 1884 42472 1915
rect 42518 1912 42524 1964
rect 42576 1952 42582 1964
rect 43901 1955 43959 1961
rect 43901 1952 43913 1955
rect 42576 1924 43913 1952
rect 42576 1912 42582 1924
rect 43901 1921 43913 1924
rect 43947 1921 43959 1955
rect 43901 1915 43959 1921
rect 47026 1912 47032 1964
rect 47084 1912 47090 1964
rect 47762 1912 47768 1964
rect 47820 1912 47826 1964
rect 47946 1912 47952 1964
rect 48004 1912 48010 1964
rect 50522 1912 50528 1964
rect 50580 1912 50586 1964
rect 50724 1961 50752 1992
rect 62117 1989 62129 2023
rect 62163 2020 62175 2023
rect 62390 2020 62396 2032
rect 62163 1992 62396 2020
rect 62163 1989 62175 1992
rect 62117 1983 62175 1989
rect 62390 1980 62396 1992
rect 62448 1980 62454 2032
rect 62574 1980 62580 2032
rect 62632 1980 62638 2032
rect 62666 1980 62672 2032
rect 62724 2020 62730 2032
rect 65978 2020 65984 2032
rect 62724 1992 65984 2020
rect 62724 1980 62730 1992
rect 65978 1980 65984 1992
rect 66036 1980 66042 2032
rect 67637 2023 67695 2029
rect 67637 1989 67649 2023
rect 67683 2020 67695 2023
rect 68002 2020 68008 2032
rect 67683 1992 68008 2020
rect 67683 1989 67695 1992
rect 67637 1983 67695 1989
rect 68002 1980 68008 1992
rect 68060 1980 68066 2032
rect 50709 1955 50767 1961
rect 50709 1921 50721 1955
rect 50755 1921 50767 1955
rect 50709 1915 50767 1921
rect 53098 1912 53104 1964
rect 53156 1952 53162 1964
rect 53469 1955 53527 1961
rect 53469 1952 53481 1955
rect 53156 1924 53481 1952
rect 53156 1912 53162 1924
rect 53469 1921 53481 1924
rect 53515 1921 53527 1955
rect 53469 1915 53527 1921
rect 54018 1912 54024 1964
rect 54076 1952 54082 1964
rect 54076 1924 55076 1952
rect 54076 1912 54082 1924
rect 40092 1856 42472 1884
rect 42889 1887 42947 1893
rect 40092 1844 40098 1856
rect 42889 1853 42901 1887
rect 42935 1853 42947 1887
rect 42889 1847 42947 1853
rect 36872 1788 37688 1816
rect 38841 1819 38899 1825
rect 36872 1776 36878 1788
rect 38841 1785 38853 1819
rect 38887 1816 38899 1819
rect 38887 1788 42380 1816
rect 38887 1785 38899 1788
rect 38841 1779 38899 1785
rect 41690 1748 41696 1760
rect 36556 1720 41696 1748
rect 41690 1708 41696 1720
rect 41748 1708 41754 1760
rect 42352 1748 42380 1788
rect 42426 1776 42432 1828
rect 42484 1816 42490 1828
rect 42904 1816 42932 1847
rect 43714 1844 43720 1896
rect 43772 1884 43778 1896
rect 44361 1887 44419 1893
rect 44361 1884 44373 1887
rect 43772 1856 44373 1884
rect 43772 1844 43778 1856
rect 44361 1853 44373 1856
rect 44407 1853 44419 1887
rect 44361 1847 44419 1853
rect 45925 1887 45983 1893
rect 45925 1853 45937 1887
rect 45971 1853 45983 1887
rect 45925 1847 45983 1853
rect 42484 1788 42932 1816
rect 42484 1776 42490 1788
rect 43254 1776 43260 1828
rect 43312 1816 43318 1828
rect 45940 1816 45968 1847
rect 46014 1844 46020 1896
rect 46072 1884 46078 1896
rect 46293 1887 46351 1893
rect 46293 1884 46305 1887
rect 46072 1856 46305 1884
rect 46072 1844 46078 1856
rect 46293 1853 46305 1856
rect 46339 1853 46351 1887
rect 46293 1847 46351 1853
rect 47854 1844 47860 1896
rect 47912 1884 47918 1896
rect 48409 1887 48467 1893
rect 48409 1884 48421 1887
rect 47912 1856 48421 1884
rect 47912 1844 47918 1856
rect 48409 1853 48421 1856
rect 48455 1853 48467 1887
rect 48409 1847 48467 1853
rect 48774 1844 48780 1896
rect 48832 1884 48838 1896
rect 49973 1887 50031 1893
rect 49973 1884 49985 1887
rect 48832 1856 49985 1884
rect 48832 1844 48838 1856
rect 49973 1853 49985 1856
rect 50019 1853 50031 1887
rect 49973 1847 50031 1853
rect 50614 1844 50620 1896
rect 50672 1884 50678 1896
rect 51169 1887 51227 1893
rect 51169 1884 51181 1887
rect 50672 1856 51181 1884
rect 50672 1844 50678 1856
rect 51169 1853 51181 1856
rect 51215 1853 51227 1887
rect 51169 1847 51227 1853
rect 51534 1844 51540 1896
rect 51592 1884 51598 1896
rect 53193 1887 53251 1893
rect 53193 1884 53205 1887
rect 51592 1856 53205 1884
rect 51592 1844 51598 1856
rect 53193 1853 53205 1856
rect 53239 1853 53251 1887
rect 53193 1847 53251 1853
rect 53374 1844 53380 1896
rect 53432 1884 53438 1896
rect 53929 1887 53987 1893
rect 53929 1884 53941 1887
rect 53432 1856 53941 1884
rect 53432 1844 53438 1856
rect 53929 1853 53941 1856
rect 53975 1853 53987 1887
rect 53929 1847 53987 1853
rect 54570 1844 54576 1896
rect 54628 1884 54634 1896
rect 54941 1887 54999 1893
rect 54941 1884 54953 1887
rect 54628 1856 54953 1884
rect 54628 1844 54634 1856
rect 54941 1853 54953 1856
rect 54987 1853 54999 1887
rect 55048 1884 55076 1924
rect 55766 1912 55772 1964
rect 55824 1912 55830 1964
rect 56229 1955 56287 1961
rect 56229 1952 56241 1955
rect 55876 1924 56241 1952
rect 55876 1884 55904 1924
rect 56229 1921 56241 1924
rect 56275 1921 56287 1955
rect 56229 1915 56287 1921
rect 57054 1912 57060 1964
rect 57112 1952 57118 1964
rect 57793 1955 57851 1961
rect 57793 1952 57805 1955
rect 57112 1924 57805 1952
rect 57112 1912 57118 1924
rect 57793 1921 57805 1924
rect 57839 1921 57851 1955
rect 57793 1915 57851 1921
rect 59998 1912 60004 1964
rect 60056 1912 60062 1964
rect 60090 1912 60096 1964
rect 60148 1952 60154 1964
rect 62942 1952 62948 1964
rect 60148 1924 62948 1952
rect 60148 1912 60154 1924
rect 62942 1912 62948 1924
rect 63000 1912 63006 1964
rect 63126 1952 63132 1964
rect 63052 1924 63132 1952
rect 55048 1856 55904 1884
rect 54941 1847 54999 1853
rect 56134 1844 56140 1896
rect 56192 1884 56198 1896
rect 56689 1887 56747 1893
rect 56689 1884 56701 1887
rect 56192 1856 56701 1884
rect 56192 1844 56198 1856
rect 56689 1853 56701 1856
rect 56735 1853 56747 1887
rect 56689 1847 56747 1853
rect 59814 1844 59820 1896
rect 59872 1884 59878 1896
rect 60737 1887 60795 1893
rect 60737 1884 60749 1887
rect 59872 1856 60749 1884
rect 59872 1844 59878 1856
rect 60737 1853 60749 1856
rect 60783 1853 60795 1887
rect 60737 1847 60795 1853
rect 61010 1844 61016 1896
rect 61068 1884 61074 1896
rect 63052 1884 63080 1924
rect 63126 1912 63132 1924
rect 63184 1912 63190 1964
rect 63494 1912 63500 1964
rect 63552 1912 63558 1964
rect 63678 1912 63684 1964
rect 63736 1912 63742 1964
rect 67269 1955 67327 1961
rect 67269 1921 67281 1955
rect 67315 1952 67327 1955
rect 67361 1955 67419 1961
rect 67361 1952 67373 1955
rect 67315 1924 67373 1952
rect 67315 1921 67327 1924
rect 67269 1915 67327 1921
rect 67361 1921 67373 1924
rect 67407 1921 67419 1955
rect 68756 1952 68784 2060
rect 69109 2057 69121 2091
rect 69155 2088 69167 2091
rect 70670 2088 70676 2100
rect 69155 2060 70676 2088
rect 69155 2057 69167 2060
rect 69109 2051 69167 2057
rect 70670 2048 70676 2060
rect 70728 2048 70734 2100
rect 69198 1980 69204 2032
rect 69256 1980 69262 2032
rect 70026 1980 70032 2032
rect 70084 2020 70090 2032
rect 71133 2023 71191 2029
rect 71133 2020 71145 2023
rect 70084 1992 71145 2020
rect 70084 1980 70090 1992
rect 71133 1989 71145 1992
rect 71179 1989 71191 2023
rect 71133 1983 71191 1989
rect 69385 1955 69443 1961
rect 69385 1952 69397 1955
rect 67361 1915 67419 1921
rect 67468 1924 68692 1952
rect 68756 1924 69397 1952
rect 61068 1856 63080 1884
rect 61068 1844 61074 1856
rect 63218 1844 63224 1896
rect 63276 1884 63282 1896
rect 64141 1887 64199 1893
rect 64141 1884 64153 1887
rect 63276 1856 64153 1884
rect 63276 1844 63282 1856
rect 64141 1853 64153 1856
rect 64187 1853 64199 1887
rect 64141 1847 64199 1853
rect 65334 1844 65340 1896
rect 65392 1884 65398 1896
rect 65705 1887 65763 1893
rect 65705 1884 65717 1887
rect 65392 1856 65717 1884
rect 65392 1844 65398 1856
rect 65705 1853 65717 1856
rect 65751 1853 65763 1887
rect 65705 1847 65763 1853
rect 66349 1887 66407 1893
rect 66349 1853 66361 1887
rect 66395 1884 66407 1887
rect 66625 1887 66683 1893
rect 66625 1884 66637 1887
rect 66395 1856 66637 1884
rect 66395 1853 66407 1856
rect 66349 1847 66407 1853
rect 66625 1853 66637 1856
rect 66671 1853 66683 1887
rect 66625 1847 66683 1853
rect 67174 1844 67180 1896
rect 67232 1884 67238 1896
rect 67468 1884 67496 1924
rect 67232 1856 67496 1884
rect 68557 1887 68615 1893
rect 67232 1844 67238 1856
rect 68557 1853 68569 1887
rect 68603 1853 68615 1887
rect 68664 1884 68692 1924
rect 69385 1921 69397 1924
rect 69431 1921 69443 1955
rect 69385 1915 69443 1921
rect 70854 1912 70860 1964
rect 70912 1912 70918 1964
rect 71406 1912 71412 1964
rect 71464 1912 71470 1964
rect 69845 1887 69903 1893
rect 69845 1884 69857 1887
rect 68664 1856 69857 1884
rect 68557 1847 68615 1853
rect 69845 1853 69857 1856
rect 69891 1853 69903 1887
rect 69845 1847 69903 1853
rect 43312 1788 45968 1816
rect 47213 1819 47271 1825
rect 43312 1776 43318 1788
rect 47213 1785 47225 1819
rect 47259 1816 47271 1819
rect 55214 1816 55220 1828
rect 47259 1788 55220 1816
rect 47259 1785 47271 1788
rect 47213 1779 47271 1785
rect 55214 1776 55220 1788
rect 55272 1776 55278 1828
rect 56045 1819 56103 1825
rect 56045 1785 56057 1819
rect 56091 1816 56103 1819
rect 62393 1819 62451 1825
rect 56091 1788 60734 1816
rect 56091 1785 56103 1788
rect 56045 1779 56103 1785
rect 51258 1748 51264 1760
rect 42352 1720 51264 1748
rect 51258 1708 51264 1720
rect 51316 1708 51322 1760
rect 58434 1708 58440 1760
rect 58492 1708 58498 1760
rect 60706 1748 60734 1788
rect 62393 1785 62405 1819
rect 62439 1816 62451 1819
rect 62439 1788 63632 1816
rect 62439 1785 62451 1788
rect 62393 1779 62451 1785
rect 63402 1748 63408 1760
rect 60706 1720 63408 1748
rect 63402 1708 63408 1720
rect 63460 1708 63466 1760
rect 63604 1748 63632 1788
rect 63770 1776 63776 1828
rect 63828 1816 63834 1828
rect 66162 1816 66168 1828
rect 63828 1788 66168 1816
rect 63828 1776 63834 1788
rect 66162 1776 66168 1788
rect 66220 1776 66226 1828
rect 68572 1816 68600 1847
rect 71314 1844 71320 1896
rect 71372 1884 71378 1896
rect 71869 1887 71927 1893
rect 71869 1884 71881 1887
rect 71372 1856 71881 1884
rect 71372 1844 71378 1856
rect 71869 1853 71881 1856
rect 71915 1853 71927 1887
rect 71869 1847 71927 1853
rect 69382 1816 69388 1828
rect 68572 1788 69388 1816
rect 69382 1776 69388 1788
rect 69440 1776 69446 1828
rect 67358 1748 67364 1760
rect 63604 1720 67364 1748
rect 67358 1708 67364 1720
rect 67416 1708 67422 1760
rect 1012 1658 74980 1680
rect 1012 1606 1858 1658
rect 1910 1606 1922 1658
rect 1974 1606 1986 1658
rect 2038 1606 2050 1658
rect 2102 1606 2114 1658
rect 2166 1606 11858 1658
rect 11910 1606 11922 1658
rect 11974 1606 11986 1658
rect 12038 1606 12050 1658
rect 12102 1606 12114 1658
rect 12166 1606 21858 1658
rect 21910 1606 21922 1658
rect 21974 1606 21986 1658
rect 22038 1606 22050 1658
rect 22102 1606 22114 1658
rect 22166 1606 31858 1658
rect 31910 1606 31922 1658
rect 31974 1606 31986 1658
rect 32038 1606 32050 1658
rect 32102 1606 32114 1658
rect 32166 1606 41858 1658
rect 41910 1606 41922 1658
rect 41974 1606 41986 1658
rect 42038 1606 42050 1658
rect 42102 1606 42114 1658
rect 42166 1606 51858 1658
rect 51910 1606 51922 1658
rect 51974 1606 51986 1658
rect 52038 1606 52050 1658
rect 52102 1606 52114 1658
rect 52166 1606 61858 1658
rect 61910 1606 61922 1658
rect 61974 1606 61986 1658
rect 62038 1606 62050 1658
rect 62102 1606 62114 1658
rect 62166 1606 71858 1658
rect 71910 1606 71922 1658
rect 71974 1606 71986 1658
rect 72038 1606 72050 1658
rect 72102 1606 72114 1658
rect 72166 1606 74980 1658
rect 1012 1584 74980 1606
rect 25406 1504 25412 1556
rect 25464 1544 25470 1556
rect 29454 1544 29460 1556
rect 25464 1516 29460 1544
rect 25464 1504 25470 1516
rect 29454 1504 29460 1516
rect 29512 1504 29518 1556
rect 30377 1547 30435 1553
rect 30377 1513 30389 1547
rect 30423 1544 30435 1547
rect 31478 1544 31484 1556
rect 30423 1516 31484 1544
rect 30423 1513 30435 1516
rect 30377 1507 30435 1513
rect 31478 1504 31484 1516
rect 31536 1504 31542 1556
rect 32858 1544 32864 1556
rect 31726 1516 32864 1544
rect 25130 1436 25136 1488
rect 25188 1476 25194 1488
rect 30466 1476 30472 1488
rect 25188 1448 30472 1476
rect 25188 1436 25194 1448
rect 30466 1436 30472 1448
rect 30524 1436 30530 1488
rect 31726 1476 31754 1516
rect 32858 1504 32864 1516
rect 32916 1504 32922 1556
rect 35437 1547 35495 1553
rect 35437 1513 35449 1547
rect 35483 1544 35495 1547
rect 35618 1544 35624 1556
rect 35483 1516 35624 1544
rect 35483 1513 35495 1516
rect 35437 1507 35495 1513
rect 35618 1504 35624 1516
rect 35676 1504 35682 1556
rect 38105 1547 38163 1553
rect 38105 1513 38117 1547
rect 38151 1544 38163 1547
rect 38746 1544 38752 1556
rect 38151 1516 38752 1544
rect 38151 1513 38163 1516
rect 38105 1507 38163 1513
rect 38746 1504 38752 1516
rect 38804 1504 38810 1556
rect 41230 1504 41236 1556
rect 41288 1504 41294 1556
rect 59078 1504 59084 1556
rect 59136 1504 59142 1556
rect 59170 1504 59176 1556
rect 59228 1544 59234 1556
rect 59228 1516 64874 1544
rect 59228 1504 59234 1516
rect 30576 1448 31754 1476
rect 23934 1368 23940 1420
rect 23992 1408 23998 1420
rect 24489 1411 24547 1417
rect 24489 1408 24501 1411
rect 23992 1380 24501 1408
rect 23992 1368 23998 1380
rect 24489 1377 24501 1380
rect 24535 1377 24547 1411
rect 30576 1408 30604 1448
rect 32674 1436 32680 1488
rect 32732 1476 32738 1488
rect 34882 1476 34888 1488
rect 32732 1448 34888 1476
rect 32732 1436 32738 1448
rect 34882 1436 34888 1448
rect 34940 1436 34946 1488
rect 47578 1436 47584 1488
rect 47636 1476 47642 1488
rect 55950 1476 55956 1488
rect 47636 1448 55956 1476
rect 47636 1436 47642 1448
rect 55950 1436 55956 1448
rect 56008 1436 56014 1488
rect 60550 1436 60556 1488
rect 60608 1436 60614 1488
rect 62117 1479 62175 1485
rect 62117 1445 62129 1479
rect 62163 1476 62175 1479
rect 62390 1476 62396 1488
rect 62163 1448 62396 1476
rect 62163 1445 62175 1448
rect 62117 1439 62175 1445
rect 62390 1436 62396 1448
rect 62448 1436 62454 1488
rect 63494 1436 63500 1488
rect 63552 1436 63558 1488
rect 64846 1476 64874 1516
rect 66530 1504 66536 1556
rect 66588 1504 66594 1556
rect 68278 1504 68284 1556
rect 68336 1504 68342 1556
rect 69198 1504 69204 1556
rect 69256 1504 69262 1556
rect 69474 1504 69480 1556
rect 69532 1544 69538 1556
rect 69569 1547 69627 1553
rect 69569 1544 69581 1547
rect 69532 1516 69581 1544
rect 69532 1504 69538 1516
rect 69569 1513 69581 1516
rect 69615 1513 69627 1547
rect 69569 1507 69627 1513
rect 67266 1476 67272 1488
rect 64846 1448 67272 1476
rect 67266 1436 67272 1448
rect 67324 1436 67330 1488
rect 24489 1371 24547 1377
rect 29288 1380 30604 1408
rect 23474 1300 23480 1352
rect 23532 1340 23538 1352
rect 23569 1343 23627 1349
rect 23569 1340 23581 1343
rect 23532 1312 23581 1340
rect 23532 1300 23538 1312
rect 23569 1309 23581 1312
rect 23615 1309 23627 1343
rect 23569 1303 23627 1309
rect 25682 1300 25688 1352
rect 25740 1300 25746 1352
rect 26145 1343 26203 1349
rect 26145 1309 26157 1343
rect 26191 1309 26203 1343
rect 26145 1303 26203 1309
rect 26697 1343 26755 1349
rect 26697 1309 26709 1343
rect 26743 1340 26755 1343
rect 26878 1340 26884 1352
rect 26743 1312 26884 1340
rect 26743 1309 26755 1312
rect 26697 1303 26755 1309
rect 26160 1272 26188 1303
rect 26878 1300 26884 1312
rect 26936 1300 26942 1352
rect 27246 1300 27252 1352
rect 27304 1300 27310 1352
rect 29288 1349 29316 1380
rect 30834 1368 30840 1420
rect 30892 1408 30898 1420
rect 33134 1408 33140 1420
rect 30892 1380 33140 1408
rect 30892 1368 30898 1380
rect 33134 1368 33140 1380
rect 33192 1368 33198 1420
rect 35360 1380 35664 1408
rect 29273 1343 29331 1349
rect 29273 1309 29285 1343
rect 29319 1309 29331 1343
rect 29273 1303 29331 1309
rect 29822 1300 29828 1352
rect 29880 1300 29886 1352
rect 30006 1300 30012 1352
rect 30064 1340 30070 1352
rect 30469 1343 30527 1349
rect 30469 1340 30481 1343
rect 30064 1312 30481 1340
rect 30064 1300 30070 1312
rect 30469 1309 30481 1312
rect 30515 1309 30527 1343
rect 32033 1343 32091 1349
rect 32033 1340 32045 1343
rect 30469 1303 30527 1309
rect 30576 1312 32045 1340
rect 28258 1272 28264 1284
rect 26160 1244 28264 1272
rect 28258 1232 28264 1244
rect 28316 1232 28322 1284
rect 28353 1275 28411 1281
rect 28353 1241 28365 1275
rect 28399 1272 28411 1275
rect 28534 1272 28540 1284
rect 28399 1244 28540 1272
rect 28399 1241 28411 1244
rect 28353 1235 28411 1241
rect 28534 1232 28540 1244
rect 28592 1232 28598 1284
rect 30576 1272 30604 1312
rect 32033 1309 32045 1312
rect 32079 1309 32091 1343
rect 32033 1303 32091 1309
rect 32677 1343 32735 1349
rect 32677 1309 32689 1343
rect 32723 1340 32735 1343
rect 32769 1343 32827 1349
rect 32769 1340 32781 1343
rect 32723 1312 32781 1340
rect 32723 1309 32735 1312
rect 32677 1303 32735 1309
rect 32769 1309 32781 1312
rect 32815 1309 32827 1343
rect 32769 1303 32827 1309
rect 33962 1300 33968 1352
rect 34020 1300 34026 1352
rect 34885 1343 34943 1349
rect 34885 1309 34897 1343
rect 34931 1340 34943 1343
rect 35360 1340 35388 1380
rect 34931 1312 35388 1340
rect 34931 1309 34943 1312
rect 34885 1303 34943 1309
rect 35434 1300 35440 1352
rect 35492 1340 35498 1352
rect 35529 1343 35587 1349
rect 35529 1340 35541 1343
rect 35492 1312 35541 1340
rect 35492 1300 35498 1312
rect 35529 1309 35541 1312
rect 35575 1309 35587 1343
rect 35636 1340 35664 1380
rect 38120 1380 38332 1408
rect 36354 1340 36360 1352
rect 35636 1312 36360 1340
rect 35529 1303 35587 1309
rect 36354 1300 36360 1312
rect 36412 1300 36418 1352
rect 37553 1343 37611 1349
rect 37553 1309 37565 1343
rect 37599 1340 37611 1343
rect 38120 1340 38148 1380
rect 37599 1312 38148 1340
rect 37599 1309 37611 1312
rect 37553 1303 37611 1309
rect 38194 1300 38200 1352
rect 38252 1300 38258 1352
rect 38304 1340 38332 1380
rect 40494 1368 40500 1420
rect 40552 1408 40558 1420
rect 41414 1408 41420 1420
rect 40552 1380 41420 1408
rect 40552 1368 40558 1380
rect 41414 1368 41420 1380
rect 41472 1368 41478 1420
rect 46661 1411 46719 1417
rect 46661 1408 46673 1411
rect 46124 1380 46673 1408
rect 38654 1340 38660 1352
rect 38304 1312 38660 1340
rect 38654 1300 38660 1312
rect 38712 1300 38718 1352
rect 39758 1300 39764 1352
rect 39816 1300 39822 1352
rect 40034 1300 40040 1352
rect 40092 1340 40098 1352
rect 41785 1343 41843 1349
rect 41785 1340 41797 1343
rect 40092 1312 41797 1340
rect 40092 1300 40098 1312
rect 41785 1309 41797 1312
rect 41831 1309 41843 1343
rect 41785 1303 41843 1309
rect 42334 1300 42340 1352
rect 42392 1300 42398 1352
rect 42702 1300 42708 1352
rect 42760 1340 42766 1352
rect 43809 1343 43867 1349
rect 43809 1340 43821 1343
rect 42760 1312 43821 1340
rect 42760 1300 42766 1312
rect 43809 1309 43821 1312
rect 43855 1309 43867 1343
rect 43809 1303 43867 1309
rect 43898 1300 43904 1352
rect 43956 1340 43962 1352
rect 44361 1343 44419 1349
rect 44361 1340 44373 1343
rect 43956 1312 44373 1340
rect 43956 1300 43962 1312
rect 44361 1309 44373 1312
rect 44407 1309 44419 1343
rect 44361 1303 44419 1309
rect 45186 1300 45192 1352
rect 45244 1300 45250 1352
rect 45462 1300 45468 1352
rect 45520 1340 45526 1352
rect 46124 1340 46152 1380
rect 46661 1377 46673 1380
rect 46707 1377 46719 1411
rect 46661 1371 46719 1377
rect 49234 1368 49240 1420
rect 49292 1408 49298 1420
rect 50525 1411 50583 1417
rect 50525 1408 50537 1411
rect 49292 1380 50537 1408
rect 49292 1368 49298 1380
rect 50525 1377 50537 1380
rect 50571 1377 50583 1411
rect 50525 1371 50583 1377
rect 58434 1368 58440 1420
rect 58492 1408 58498 1420
rect 58492 1380 59400 1408
rect 58492 1368 58498 1380
rect 47213 1343 47271 1349
rect 47213 1340 47225 1343
rect 45520 1312 46152 1340
rect 46216 1312 47225 1340
rect 45520 1300 45526 1312
rect 30300 1244 30604 1272
rect 31665 1275 31723 1281
rect 23753 1207 23811 1213
rect 23753 1173 23765 1207
rect 23799 1204 23811 1207
rect 27614 1204 27620 1216
rect 23799 1176 27620 1204
rect 23799 1173 23811 1176
rect 23753 1167 23811 1173
rect 27614 1164 27620 1176
rect 27672 1164 27678 1216
rect 27801 1207 27859 1213
rect 27801 1173 27813 1207
rect 27847 1204 27859 1207
rect 30300 1204 30328 1244
rect 31665 1241 31677 1275
rect 31711 1241 31723 1275
rect 31665 1235 31723 1241
rect 27847 1176 30328 1204
rect 31680 1204 31708 1235
rect 35618 1232 35624 1284
rect 35676 1272 35682 1284
rect 36449 1275 36507 1281
rect 36449 1272 36461 1275
rect 35676 1244 36461 1272
rect 35676 1232 35682 1244
rect 36449 1241 36461 1244
rect 36495 1241 36507 1275
rect 36449 1235 36507 1241
rect 38286 1232 38292 1284
rect 38344 1272 38350 1284
rect 39117 1275 39175 1281
rect 39117 1272 39129 1275
rect 38344 1244 39129 1272
rect 38344 1232 38350 1244
rect 39117 1241 39129 1244
rect 39163 1241 39175 1275
rect 39117 1235 39175 1241
rect 39574 1232 39580 1284
rect 39632 1272 39638 1284
rect 40681 1275 40739 1281
rect 40681 1272 40693 1275
rect 39632 1244 40693 1272
rect 39632 1232 39638 1244
rect 40681 1241 40693 1244
rect 40727 1241 40739 1275
rect 40681 1235 40739 1241
rect 40954 1232 40960 1284
rect 41012 1272 41018 1284
rect 43257 1275 43315 1281
rect 43257 1272 43269 1275
rect 41012 1244 43269 1272
rect 41012 1232 41018 1244
rect 43257 1241 43269 1244
rect 43303 1241 43315 1275
rect 43257 1235 43315 1241
rect 45094 1232 45100 1284
rect 45152 1272 45158 1284
rect 46109 1275 46167 1281
rect 46109 1272 46121 1275
rect 45152 1244 46121 1272
rect 45152 1232 45158 1244
rect 46109 1241 46121 1244
rect 46155 1241 46167 1275
rect 46109 1235 46167 1241
rect 44082 1204 44088 1216
rect 31680 1176 44088 1204
rect 27847 1173 27859 1176
rect 27801 1167 27859 1173
rect 44082 1164 44088 1176
rect 44140 1164 44146 1216
rect 44634 1164 44640 1216
rect 44692 1204 44698 1216
rect 46216 1204 46244 1312
rect 47213 1309 47225 1312
rect 47259 1309 47271 1343
rect 47213 1303 47271 1309
rect 47486 1300 47492 1352
rect 47544 1300 47550 1352
rect 47762 1300 47768 1352
rect 47820 1340 47826 1352
rect 48961 1343 49019 1349
rect 48961 1340 48973 1343
rect 47820 1312 48973 1340
rect 47820 1300 47826 1312
rect 48961 1309 48973 1312
rect 49007 1309 49019 1343
rect 49513 1343 49571 1349
rect 49513 1340 49525 1343
rect 48961 1303 49019 1309
rect 49068 1312 49525 1340
rect 46474 1232 46480 1284
rect 46532 1272 46538 1284
rect 48409 1275 48467 1281
rect 48409 1272 48421 1275
rect 46532 1244 48421 1272
rect 46532 1232 46538 1244
rect 48409 1241 48421 1244
rect 48455 1241 48467 1275
rect 48409 1235 48467 1241
rect 44692 1176 46244 1204
rect 44692 1164 44698 1176
rect 48130 1164 48136 1216
rect 48188 1204 48194 1216
rect 49068 1204 49096 1312
rect 49513 1309 49525 1312
rect 49559 1309 49571 1343
rect 49513 1303 49571 1309
rect 49602 1300 49608 1352
rect 49660 1340 49666 1352
rect 50065 1343 50123 1349
rect 50065 1340 50077 1343
rect 49660 1312 50077 1340
rect 49660 1300 49666 1312
rect 50065 1309 50077 1312
rect 50111 1309 50123 1343
rect 50065 1303 50123 1309
rect 50798 1300 50804 1352
rect 50856 1340 50862 1352
rect 52089 1343 52147 1349
rect 52089 1340 52101 1343
rect 50856 1312 52101 1340
rect 50856 1300 50862 1312
rect 52089 1309 52101 1312
rect 52135 1309 52147 1343
rect 52089 1303 52147 1309
rect 52270 1300 52276 1352
rect 52328 1340 52334 1352
rect 52641 1343 52699 1349
rect 52641 1340 52653 1343
rect 52328 1312 52653 1340
rect 52328 1300 52334 1312
rect 52641 1309 52653 1312
rect 52687 1309 52699 1343
rect 52641 1303 52699 1309
rect 53650 1300 53656 1352
rect 53708 1340 53714 1352
rect 54113 1343 54171 1349
rect 54113 1340 54125 1343
rect 53708 1312 54125 1340
rect 53708 1300 53714 1312
rect 54113 1309 54125 1312
rect 54159 1309 54171 1343
rect 54113 1303 54171 1309
rect 54665 1343 54723 1349
rect 54665 1309 54677 1343
rect 54711 1309 54723 1343
rect 54665 1303 54723 1309
rect 49142 1232 49148 1284
rect 49200 1272 49206 1284
rect 51718 1272 51724 1284
rect 49200 1244 51724 1272
rect 49200 1232 49206 1244
rect 51718 1232 51724 1244
rect 51776 1232 51782 1284
rect 52362 1232 52368 1284
rect 52420 1272 52426 1284
rect 53561 1275 53619 1281
rect 53561 1272 53573 1275
rect 52420 1244 53573 1272
rect 52420 1232 52426 1244
rect 53561 1241 53573 1244
rect 53607 1241 53619 1275
rect 53561 1235 53619 1241
rect 48188 1176 49096 1204
rect 48188 1164 48194 1176
rect 50522 1164 50528 1216
rect 50580 1204 50586 1216
rect 51537 1207 51595 1213
rect 51537 1204 51549 1207
rect 50580 1176 51549 1204
rect 50580 1164 50586 1176
rect 51537 1173 51549 1176
rect 51583 1173 51595 1207
rect 51537 1167 51595 1173
rect 52914 1164 52920 1216
rect 52972 1204 52978 1216
rect 54680 1204 54708 1303
rect 54846 1300 54852 1352
rect 54904 1340 54910 1352
rect 55217 1343 55275 1349
rect 55217 1340 55229 1343
rect 54904 1312 55229 1340
rect 54904 1300 54910 1312
rect 55217 1309 55229 1312
rect 55263 1309 55275 1343
rect 55217 1303 55275 1309
rect 56318 1300 56324 1352
rect 56376 1340 56382 1352
rect 56689 1343 56747 1349
rect 56689 1340 56701 1343
rect 56376 1312 56701 1340
rect 56376 1300 56382 1312
rect 56689 1309 56701 1312
rect 56735 1309 56747 1343
rect 56689 1303 56747 1309
rect 57241 1343 57299 1349
rect 57241 1309 57253 1343
rect 57287 1309 57299 1343
rect 57241 1303 57299 1309
rect 54754 1232 54760 1284
rect 54812 1272 54818 1284
rect 56137 1275 56195 1281
rect 56137 1272 56149 1275
rect 54812 1244 56149 1272
rect 54812 1232 54818 1244
rect 56137 1241 56149 1244
rect 56183 1241 56195 1275
rect 56137 1235 56195 1241
rect 52972 1176 54708 1204
rect 52972 1164 52978 1176
rect 55674 1164 55680 1216
rect 55732 1204 55738 1216
rect 57256 1204 57284 1303
rect 59262 1300 59268 1352
rect 59320 1300 59326 1352
rect 59372 1340 59400 1380
rect 63604 1380 63816 1408
rect 59817 1343 59875 1349
rect 59817 1340 59829 1343
rect 59372 1312 59829 1340
rect 59817 1309 59829 1312
rect 59863 1309 59875 1343
rect 59817 1303 59875 1309
rect 61194 1300 61200 1352
rect 61252 1340 61258 1352
rect 61289 1343 61347 1349
rect 61289 1340 61301 1343
rect 61252 1312 61301 1340
rect 61252 1300 61258 1312
rect 61289 1309 61301 1312
rect 61335 1309 61347 1343
rect 61289 1303 61347 1309
rect 61933 1343 61991 1349
rect 61933 1309 61945 1343
rect 61979 1340 61991 1343
rect 62298 1340 62304 1352
rect 61979 1312 62304 1340
rect 61979 1309 61991 1312
rect 61933 1303 61991 1309
rect 62298 1300 62304 1312
rect 62356 1300 62362 1352
rect 62574 1300 62580 1352
rect 62632 1340 62638 1352
rect 63604 1340 63632 1380
rect 62632 1312 63632 1340
rect 62632 1300 62638 1312
rect 63678 1300 63684 1352
rect 63736 1300 63742 1352
rect 63788 1340 63816 1380
rect 69934 1368 69940 1420
rect 69992 1408 69998 1420
rect 71133 1411 71191 1417
rect 71133 1408 71145 1411
rect 69992 1380 71145 1408
rect 69992 1368 69998 1380
rect 71133 1377 71145 1380
rect 71179 1377 71191 1411
rect 71133 1371 71191 1377
rect 66073 1343 66131 1349
rect 66073 1340 66085 1343
rect 63788 1312 66085 1340
rect 66073 1309 66085 1312
rect 66119 1309 66131 1343
rect 66073 1303 66131 1309
rect 66714 1300 66720 1352
rect 66772 1340 66778 1352
rect 66993 1343 67051 1349
rect 66993 1340 67005 1343
rect 66772 1312 67005 1340
rect 66772 1300 66778 1312
rect 66993 1309 67005 1312
rect 67039 1309 67051 1343
rect 66993 1303 67051 1309
rect 67634 1300 67640 1352
rect 67692 1300 67698 1352
rect 68094 1300 68100 1352
rect 68152 1340 68158 1352
rect 70121 1343 70179 1349
rect 70121 1340 70133 1343
rect 68152 1312 70133 1340
rect 68152 1300 68158 1312
rect 70121 1309 70133 1312
rect 70167 1309 70179 1343
rect 70121 1303 70179 1309
rect 70578 1300 70584 1352
rect 70636 1340 70642 1352
rect 70673 1343 70731 1349
rect 70673 1340 70685 1343
rect 70636 1312 70685 1340
rect 70636 1300 70642 1312
rect 70673 1309 70685 1312
rect 70719 1309 70731 1343
rect 70673 1303 70731 1309
rect 70854 1300 70860 1352
rect 70912 1340 70918 1352
rect 72145 1343 72203 1349
rect 72145 1340 72157 1343
rect 70912 1312 72157 1340
rect 70912 1300 70918 1312
rect 72145 1309 72157 1312
rect 72191 1309 72203 1343
rect 72145 1303 72203 1309
rect 72789 1343 72847 1349
rect 72789 1309 72801 1343
rect 72835 1340 72847 1343
rect 73801 1343 73859 1349
rect 73801 1340 73813 1343
rect 72835 1312 73813 1340
rect 72835 1309 72847 1312
rect 72789 1303 72847 1309
rect 73801 1309 73813 1312
rect 73847 1309 73859 1343
rect 73801 1303 73859 1309
rect 64598 1232 64604 1284
rect 64656 1232 64662 1284
rect 65426 1232 65432 1284
rect 65484 1272 65490 1284
rect 65521 1275 65579 1281
rect 65521 1272 65533 1275
rect 65484 1244 65533 1272
rect 65484 1232 65490 1244
rect 65521 1241 65533 1244
rect 65567 1241 65579 1275
rect 65521 1235 65579 1241
rect 67542 1232 67548 1284
rect 67600 1272 67606 1284
rect 68189 1275 68247 1281
rect 68189 1272 68201 1275
rect 67600 1244 68201 1272
rect 67600 1232 67606 1244
rect 68189 1241 68201 1244
rect 68235 1241 68247 1275
rect 68189 1235 68247 1241
rect 72602 1232 72608 1284
rect 72660 1272 72666 1284
rect 73249 1275 73307 1281
rect 73249 1272 73261 1275
rect 72660 1244 73261 1272
rect 72660 1232 72666 1244
rect 73249 1241 73261 1244
rect 73295 1241 73307 1275
rect 73249 1235 73307 1241
rect 55732 1176 57284 1204
rect 55732 1164 55738 1176
rect 57330 1164 57336 1216
rect 57388 1204 57394 1216
rect 65610 1204 65616 1216
rect 57388 1176 65616 1204
rect 57388 1164 57394 1176
rect 65610 1164 65616 1176
rect 65668 1164 65674 1216
rect 1012 1114 74980 1136
rect 1012 1062 4210 1114
rect 4262 1062 4274 1114
rect 4326 1062 4338 1114
rect 4390 1062 4402 1114
rect 4454 1062 4466 1114
rect 4518 1062 14210 1114
rect 14262 1062 14274 1114
rect 14326 1062 14338 1114
rect 14390 1062 14402 1114
rect 14454 1062 14466 1114
rect 14518 1062 24210 1114
rect 24262 1062 24274 1114
rect 24326 1062 24338 1114
rect 24390 1062 24402 1114
rect 24454 1062 24466 1114
rect 24518 1062 34210 1114
rect 34262 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 44210 1114
rect 44262 1062 44274 1114
rect 44326 1062 44338 1114
rect 44390 1062 44402 1114
rect 44454 1062 44466 1114
rect 44518 1062 54210 1114
rect 54262 1062 54274 1114
rect 54326 1062 54338 1114
rect 54390 1062 54402 1114
rect 54454 1062 54466 1114
rect 54518 1062 64210 1114
rect 64262 1062 64274 1114
rect 64326 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 74210 1114
rect 74262 1062 74274 1114
rect 74326 1062 74338 1114
rect 74390 1062 74402 1114
rect 74454 1062 74466 1114
rect 74518 1062 74980 1114
rect 1012 1040 74980 1062
rect 25682 960 25688 1012
rect 25740 1000 25746 1012
rect 25740 972 26234 1000
rect 25740 960 25746 972
rect 26206 796 26234 972
rect 28258 960 28264 1012
rect 28316 1000 28322 1012
rect 30834 1000 30840 1012
rect 28316 972 30840 1000
rect 28316 960 28322 972
rect 30834 960 30840 972
rect 30892 960 30898 1012
rect 33318 960 33324 1012
rect 33376 1000 33382 1012
rect 33376 972 34652 1000
rect 33376 960 33382 972
rect 29822 892 29828 944
rect 29880 932 29886 944
rect 34514 932 34520 944
rect 29880 904 34520 932
rect 29880 892 29886 904
rect 34514 892 34520 904
rect 34572 892 34578 944
rect 34624 932 34652 972
rect 41414 960 41420 1012
rect 41472 1000 41478 1012
rect 43898 1000 43904 1012
rect 41472 972 43904 1000
rect 41472 960 41478 972
rect 43898 960 43904 972
rect 43956 960 43962 1012
rect 44082 960 44088 1012
rect 44140 1000 44146 1012
rect 49142 1000 49148 1012
rect 44140 972 49148 1000
rect 44140 960 44146 972
rect 49142 960 49148 972
rect 49200 960 49206 1012
rect 51718 960 51724 1012
rect 51776 1000 51782 1012
rect 57330 1000 57336 1012
rect 51776 972 57336 1000
rect 51776 960 51782 972
rect 57330 960 57336 972
rect 57388 960 57394 1012
rect 60274 960 60280 1012
rect 60332 1000 60338 1012
rect 64598 1000 64604 1012
rect 60332 972 64604 1000
rect 60332 960 60338 972
rect 64598 960 64604 972
rect 64656 960 64662 1012
rect 45186 932 45192 944
rect 34624 904 45192 932
rect 45186 892 45192 904
rect 45244 892 45250 944
rect 48498 892 48504 944
rect 48556 932 48562 944
rect 49602 932 49608 944
rect 48556 904 49608 932
rect 48556 892 48562 904
rect 49602 892 49608 904
rect 49660 892 49666 944
rect 27246 824 27252 876
rect 27304 864 27310 876
rect 32582 864 32588 876
rect 27304 836 32588 864
rect 27304 824 27310 836
rect 32582 824 32588 836
rect 32640 824 32646 876
rect 47486 864 47492 876
rect 38626 836 47492 864
rect 33410 796 33416 808
rect 26206 768 33416 796
rect 33410 756 33416 768
rect 33468 756 33474 808
rect 30926 688 30932 740
rect 30984 728 30990 740
rect 38626 728 38654 836
rect 47486 824 47492 836
rect 47544 824 47550 876
rect 30984 700 38654 728
rect 30984 688 30990 700
rect 23106 76 23112 128
rect 23164 116 23170 128
rect 65702 116 65708 128
rect 23164 88 65708 116
rect 23164 76 23170 88
rect 65702 76 65708 88
rect 65760 76 65766 128
<< via1 >>
rect 74210 85926 74262 85978
rect 74274 85926 74326 85978
rect 74338 85926 74390 85978
rect 74402 85926 74454 85978
rect 74466 85926 74518 85978
rect 71858 85382 71910 85434
rect 71922 85382 71974 85434
rect 71986 85382 72038 85434
rect 72050 85382 72102 85434
rect 72114 85382 72166 85434
rect 74210 84838 74262 84890
rect 74274 84838 74326 84890
rect 74338 84838 74390 84890
rect 74402 84838 74454 84890
rect 74466 84838 74518 84890
rect 71858 84294 71910 84346
rect 71922 84294 71974 84346
rect 71986 84294 72038 84346
rect 72050 84294 72102 84346
rect 72114 84294 72166 84346
rect 63500 84192 63552 84244
rect 74210 83750 74262 83802
rect 74274 83750 74326 83802
rect 74338 83750 74390 83802
rect 74402 83750 74454 83802
rect 74466 83750 74518 83802
rect 71858 83206 71910 83258
rect 71922 83206 71974 83258
rect 71986 83206 72038 83258
rect 72050 83206 72102 83258
rect 72114 83206 72166 83258
rect 66904 83104 66956 83156
rect 69204 83036 69256 83088
rect 74210 82662 74262 82714
rect 74274 82662 74326 82714
rect 74338 82662 74390 82714
rect 74402 82662 74454 82714
rect 74466 82662 74518 82714
rect 63500 82356 63552 82408
rect 71858 82118 71910 82170
rect 71922 82118 71974 82170
rect 71986 82118 72038 82170
rect 72050 82118 72102 82170
rect 72114 82118 72166 82170
rect 74210 81574 74262 81626
rect 74274 81574 74326 81626
rect 74338 81574 74390 81626
rect 74402 81574 74454 81626
rect 74466 81574 74518 81626
rect 71858 81030 71910 81082
rect 71922 81030 71974 81082
rect 71986 81030 72038 81082
rect 72050 81030 72102 81082
rect 72114 81030 72166 81082
rect 66720 80928 66772 80980
rect 66996 80588 67048 80640
rect 74210 80486 74262 80538
rect 74274 80486 74326 80538
rect 74338 80486 74390 80538
rect 74402 80486 74454 80538
rect 74466 80486 74518 80538
rect 63500 79976 63552 80028
rect 71858 79942 71910 79994
rect 71922 79942 71974 79994
rect 71986 79942 72038 79994
rect 72050 79942 72102 79994
rect 72114 79942 72166 79994
rect 74210 79398 74262 79450
rect 74274 79398 74326 79450
rect 74338 79398 74390 79450
rect 74402 79398 74454 79450
rect 74466 79398 74518 79450
rect 71858 78854 71910 78906
rect 71922 78854 71974 78906
rect 71986 78854 72038 78906
rect 72050 78854 72102 78906
rect 72114 78854 72166 78906
rect 65616 78684 65668 78736
rect 67088 78412 67140 78464
rect 74210 78310 74262 78362
rect 74274 78310 74326 78362
rect 74338 78310 74390 78362
rect 74402 78310 74454 78362
rect 74466 78310 74518 78362
rect 63500 78004 63552 78056
rect 71858 77766 71910 77818
rect 71922 77766 71974 77818
rect 71986 77766 72038 77818
rect 72050 77766 72102 77818
rect 72114 77766 72166 77818
rect 63592 77392 63644 77444
rect 74210 77222 74262 77274
rect 74274 77222 74326 77274
rect 74338 77222 74390 77274
rect 74402 77222 74454 77274
rect 74466 77222 74518 77274
rect 63500 76690 63552 76742
rect 71858 76678 71910 76730
rect 71922 76678 71974 76730
rect 71986 76678 72038 76730
rect 72050 76678 72102 76730
rect 72114 76678 72166 76730
rect 63684 76100 63736 76152
rect 74210 76134 74262 76186
rect 74274 76134 74326 76186
rect 74338 76134 74390 76186
rect 74402 76134 74454 76186
rect 74466 76134 74518 76186
rect 63592 75760 63644 75812
rect 71858 75590 71910 75642
rect 71922 75590 71974 75642
rect 71986 75590 72038 75642
rect 72050 75590 72102 75642
rect 72114 75590 72166 75642
rect 74210 75046 74262 75098
rect 74274 75046 74326 75098
rect 74338 75046 74390 75098
rect 74402 75046 74454 75098
rect 74466 75046 74518 75098
rect 63868 74536 63920 74588
rect 71858 74502 71910 74554
rect 71922 74502 71974 74554
rect 71986 74502 72038 74554
rect 72050 74502 72102 74554
rect 72114 74502 72166 74554
rect 64144 73924 64196 73976
rect 74210 73958 74262 74010
rect 74274 73958 74326 74010
rect 74338 73958 74390 74010
rect 74402 73958 74454 74010
rect 74466 73958 74518 74010
rect 71858 73414 71910 73466
rect 71922 73414 71974 73466
rect 71986 73414 72038 73466
rect 72050 73414 72102 73466
rect 72114 73414 72166 73466
rect 63592 73176 63644 73228
rect 74210 72870 74262 72922
rect 74274 72870 74326 72922
rect 74338 72870 74390 72922
rect 74402 72870 74454 72922
rect 74466 72870 74518 72922
rect 71858 72326 71910 72378
rect 71922 72326 71974 72378
rect 71986 72326 72038 72378
rect 72050 72326 72102 72378
rect 72114 72326 72166 72378
rect 65708 72156 65760 72208
rect 69020 72088 69072 72140
rect 74210 71782 74262 71834
rect 74274 71782 74326 71834
rect 74338 71782 74390 71834
rect 74402 71782 74454 71834
rect 74466 71782 74518 71834
rect 63500 71612 63552 71664
rect 66168 71612 66220 71664
rect 65616 71544 65668 71596
rect 66352 71544 66404 71596
rect 63592 71408 63644 71460
rect 71858 71238 71910 71290
rect 71922 71238 71974 71290
rect 71986 71238 72038 71290
rect 72050 71238 72102 71290
rect 72114 71238 72166 71290
rect 63500 70796 63552 70848
rect 74210 70694 74262 70746
rect 74274 70694 74326 70746
rect 74338 70694 74390 70746
rect 74402 70694 74454 70746
rect 74466 70694 74518 70746
rect 71858 70150 71910 70202
rect 71922 70150 71974 70202
rect 71986 70150 72038 70202
rect 72050 70150 72102 70202
rect 72114 70150 72166 70202
rect 65616 69980 65668 70032
rect 63776 69572 63828 69624
rect 74210 69606 74262 69658
rect 74274 69606 74326 69658
rect 74338 69606 74390 69658
rect 74402 69606 74454 69658
rect 74466 69606 74518 69658
rect 71858 69062 71910 69114
rect 71922 69062 71974 69114
rect 71986 69062 72038 69114
rect 72050 69062 72102 69114
rect 72114 69062 72166 69114
rect 63500 68960 63552 69012
rect 66628 68620 66680 68672
rect 74210 68518 74262 68570
rect 74274 68518 74326 68570
rect 74338 68518 74390 68570
rect 74402 68518 74454 68570
rect 74466 68518 74518 68570
rect 71858 67974 71910 68026
rect 71922 67974 71974 68026
rect 71986 67974 72038 68026
rect 72050 67974 72102 68026
rect 72114 67974 72166 68026
rect 64788 67600 64840 67652
rect 65432 67532 65484 67584
rect 74210 67430 74262 67482
rect 74274 67430 74326 67482
rect 74338 67430 74390 67482
rect 74402 67430 74454 67482
rect 74466 67430 74518 67482
rect 71858 66886 71910 66938
rect 71922 66886 71974 66938
rect 71986 66886 72038 66938
rect 72050 66886 72102 66938
rect 72114 66886 72166 66938
rect 63592 66444 63644 66496
rect 74210 66342 74262 66394
rect 74274 66342 74326 66394
rect 74338 66342 74390 66394
rect 74402 66342 74454 66394
rect 74466 66342 74518 66394
rect 71858 65798 71910 65850
rect 71922 65798 71974 65850
rect 71986 65798 72038 65850
rect 72050 65798 72102 65850
rect 72114 65798 72166 65850
rect 65340 65628 65392 65680
rect 66996 65492 67048 65544
rect 68100 65492 68152 65544
rect 63500 65220 63552 65272
rect 74210 65254 74262 65306
rect 74274 65254 74326 65306
rect 74338 65254 74390 65306
rect 74402 65254 74454 65306
rect 74466 65254 74518 65306
rect 63592 64812 63644 64864
rect 63592 64676 63644 64728
rect 63776 64676 63828 64728
rect 71858 64710 71910 64762
rect 71922 64710 71974 64762
rect 71986 64710 72038 64762
rect 72050 64710 72102 64762
rect 72114 64710 72166 64762
rect 63776 64268 63828 64320
rect 74210 64166 74262 64218
rect 74274 64166 74326 64218
rect 74338 64166 74390 64218
rect 74402 64166 74454 64218
rect 74466 64166 74518 64218
rect 63960 63588 64012 63640
rect 71858 63622 71910 63674
rect 71922 63622 71974 63674
rect 71986 63622 72038 63674
rect 72050 63622 72102 63674
rect 72114 63622 72166 63674
rect 63500 63180 63552 63232
rect 74210 63078 74262 63130
rect 74274 63078 74326 63130
rect 74338 63078 74390 63130
rect 74402 63078 74454 63130
rect 74466 63078 74518 63130
rect 71858 62534 71910 62586
rect 71922 62534 71974 62586
rect 71986 62534 72038 62586
rect 72050 62534 72102 62586
rect 72114 62534 72166 62586
rect 63776 62092 63828 62144
rect 63960 62024 64012 62076
rect 65248 62024 65300 62076
rect 74210 61990 74262 62042
rect 74274 61990 74326 62042
rect 74338 61990 74390 62042
rect 74402 61990 74454 62042
rect 74466 61990 74518 62042
rect 71858 61446 71910 61498
rect 71922 61446 71974 61498
rect 71986 61446 72038 61498
rect 72050 61446 72102 61498
rect 72114 61446 72166 61498
rect 63960 61276 64012 61328
rect 63500 61004 63552 61056
rect 74210 60902 74262 60954
rect 74274 60902 74326 60954
rect 74338 60902 74390 60954
rect 74402 60902 74454 60954
rect 74466 60902 74518 60954
rect 71858 60358 71910 60410
rect 71922 60358 71974 60410
rect 71986 60358 72038 60410
rect 72050 60358 72102 60410
rect 72114 60358 72166 60410
rect 63776 59916 63828 59968
rect 74210 59814 74262 59866
rect 74274 59814 74326 59866
rect 74338 59814 74390 59866
rect 74402 59814 74454 59866
rect 74466 59814 74518 59866
rect 71858 59270 71910 59322
rect 71922 59270 71974 59322
rect 71986 59270 72038 59322
rect 72050 59270 72102 59322
rect 72114 59270 72166 59322
rect 65156 59100 65208 59152
rect 63500 58692 63552 58744
rect 74210 58726 74262 58778
rect 74274 58726 74326 58778
rect 74338 58726 74390 58778
rect 74402 58726 74454 58778
rect 74466 58726 74518 58778
rect 71858 58182 71910 58234
rect 71922 58182 71974 58234
rect 71986 58182 72038 58234
rect 72050 58182 72102 58234
rect 72114 58182 72166 58234
rect 63776 57944 63828 57996
rect 74210 57638 74262 57690
rect 74274 57638 74326 57690
rect 74338 57638 74390 57690
rect 74402 57638 74454 57690
rect 74466 57638 74518 57690
rect 71858 57094 71910 57146
rect 71922 57094 71974 57146
rect 71986 57094 72038 57146
rect 72050 57094 72102 57146
rect 72114 57094 72166 57146
rect 65064 56924 65116 56976
rect 63500 56652 63552 56704
rect 74210 56550 74262 56602
rect 74274 56550 74326 56602
rect 74338 56550 74390 56602
rect 74402 56550 74454 56602
rect 74466 56550 74518 56602
rect 71858 56006 71910 56058
rect 71922 56006 71974 56058
rect 71986 56006 72038 56058
rect 72050 56006 72102 56058
rect 72114 56006 72166 56058
rect 63776 55564 63828 55616
rect 74210 55462 74262 55514
rect 74274 55462 74326 55514
rect 74338 55462 74390 55514
rect 74402 55462 74454 55514
rect 74466 55462 74518 55514
rect 63960 55224 64012 55276
rect 64972 55224 65024 55276
rect 71858 54918 71910 54970
rect 71922 54918 71974 54970
rect 71986 54918 72038 54970
rect 72050 54918 72102 54970
rect 72114 54918 72166 54970
rect 64052 54748 64104 54800
rect 63500 54612 63552 54664
rect 74210 54374 74262 54426
rect 74274 54374 74326 54426
rect 74338 54374 74390 54426
rect 74402 54374 74454 54426
rect 74466 54374 74518 54426
rect 71858 53830 71910 53882
rect 71922 53830 71974 53882
rect 71986 53830 72038 53882
rect 72050 53830 72102 53882
rect 72114 53830 72166 53882
rect 63776 53524 63828 53576
rect 74210 53286 74262 53338
rect 74274 53286 74326 53338
rect 74338 53286 74390 53338
rect 74402 53286 74454 53338
rect 74466 53286 74518 53338
rect 66996 53116 67048 53168
rect 71858 52742 71910 52794
rect 71922 52742 71974 52794
rect 71986 52742 72038 52794
rect 72050 52742 72102 52794
rect 72114 52742 72166 52794
rect 64696 52640 64748 52692
rect 63500 52572 63552 52624
rect 69296 52572 69348 52624
rect 74210 52198 74262 52250
rect 74274 52198 74326 52250
rect 74338 52198 74390 52250
rect 74402 52198 74454 52250
rect 74466 52198 74518 52250
rect 63500 52068 63552 52120
rect 71858 51654 71910 51706
rect 71922 51654 71974 51706
rect 71986 51654 72038 51706
rect 72050 51654 72102 51706
rect 72114 51654 72166 51706
rect 63776 51484 63828 51536
rect 66536 51484 66588 51536
rect 74210 51110 74262 51162
rect 74274 51110 74326 51162
rect 74338 51110 74390 51162
rect 74402 51110 74454 51162
rect 74466 51110 74518 51162
rect 71858 50566 71910 50618
rect 71922 50566 71974 50618
rect 71986 50566 72038 50618
rect 72050 50566 72102 50618
rect 72114 50566 72166 50618
rect 64880 50396 64932 50448
rect 69112 50328 69164 50380
rect 74210 50022 74262 50074
rect 74274 50022 74326 50074
rect 74338 50022 74390 50074
rect 74402 50022 74454 50074
rect 74466 50022 74518 50074
rect 71858 49478 71910 49530
rect 71922 49478 71974 49530
rect 71986 49478 72038 49530
rect 72050 49478 72102 49530
rect 72114 49478 72166 49530
rect 64328 48764 64380 48816
rect 74210 48934 74262 48986
rect 74274 48934 74326 48986
rect 74338 48934 74390 48986
rect 74402 48934 74454 48986
rect 74466 48934 74518 48986
rect 71858 48390 71910 48442
rect 71922 48390 71974 48442
rect 71986 48390 72038 48442
rect 72050 48390 72102 48442
rect 72114 48390 72166 48442
rect 68560 48084 68612 48136
rect 74210 47846 74262 47898
rect 74274 47846 74326 47898
rect 74338 47846 74390 47898
rect 74402 47846 74454 47898
rect 74466 47846 74518 47898
rect 64420 47676 64472 47728
rect 65524 47472 65576 47524
rect 71858 47302 71910 47354
rect 71922 47302 71974 47354
rect 71986 47302 72038 47354
rect 72050 47302 72102 47354
rect 72114 47302 72166 47354
rect 66076 47064 66128 47116
rect 65708 47039 65760 47048
rect 65708 47005 65717 47039
rect 65717 47005 65751 47039
rect 65751 47005 65760 47039
rect 65708 46996 65760 47005
rect 65984 47039 66036 47048
rect 65984 47005 65993 47039
rect 65993 47005 66027 47039
rect 66027 47005 66036 47039
rect 65984 46996 66036 47005
rect 74210 46758 74262 46810
rect 74274 46758 74326 46810
rect 74338 46758 74390 46810
rect 74402 46758 74454 46810
rect 74466 46758 74518 46810
rect 71858 46214 71910 46266
rect 71922 46214 71974 46266
rect 71986 46214 72038 46266
rect 72050 46214 72102 46266
rect 72114 46214 72166 46266
rect 65800 45908 65852 45960
rect 74210 45670 74262 45722
rect 74274 45670 74326 45722
rect 74338 45670 74390 45722
rect 74402 45670 74454 45722
rect 74466 45670 74518 45722
rect 65984 45568 66036 45620
rect 66444 45228 66496 45280
rect 71858 45126 71910 45178
rect 71922 45126 71974 45178
rect 71986 45126 72038 45178
rect 72050 45126 72102 45178
rect 72114 45126 72166 45178
rect 67180 44820 67232 44872
rect 63684 44684 63736 44736
rect 64236 44684 64288 44736
rect 63684 44548 63736 44600
rect 74210 44582 74262 44634
rect 74274 44582 74326 44634
rect 74338 44582 74390 44634
rect 74402 44582 74454 44634
rect 74466 44582 74518 44634
rect 67548 44140 67600 44192
rect 71858 44038 71910 44090
rect 71922 44038 71974 44090
rect 71986 44038 72038 44090
rect 72050 44038 72102 44090
rect 72114 44038 72166 44090
rect 64604 43800 64656 43852
rect 65524 43596 65576 43648
rect 65892 43596 65944 43648
rect 74210 43494 74262 43546
rect 74274 43494 74326 43546
rect 74338 43494 74390 43546
rect 74402 43494 74454 43546
rect 74466 43494 74518 43546
rect 64052 43392 64104 43444
rect 65524 43392 65576 43444
rect 69388 43256 69440 43308
rect 71858 42950 71910 43002
rect 71922 42950 71974 43002
rect 71986 42950 72038 43002
rect 72050 42950 72102 43002
rect 72114 42950 72166 43002
rect 63776 42780 63828 42832
rect 66904 42712 66956 42764
rect 69664 42644 69716 42696
rect 74210 42406 74262 42458
rect 74274 42406 74326 42458
rect 74338 42406 74390 42458
rect 74402 42406 74454 42458
rect 74466 42406 74518 42458
rect 71858 41862 71910 41914
rect 71922 41862 71974 41914
rect 71986 41862 72038 41914
rect 72050 41862 72102 41914
rect 72114 41862 72166 41914
rect 66720 41803 66772 41812
rect 66720 41769 66729 41803
rect 66729 41769 66763 41803
rect 66763 41769 66772 41803
rect 66720 41760 66772 41769
rect 63500 41692 63552 41744
rect 69848 41556 69900 41608
rect 74210 41318 74262 41370
rect 74274 41318 74326 41370
rect 74338 41318 74390 41370
rect 74402 41318 74454 41370
rect 74466 41318 74518 41370
rect 63960 40944 64012 40996
rect 65892 40876 65944 40928
rect 66260 40876 66312 40928
rect 71858 40774 71910 40826
rect 71922 40774 71974 40826
rect 71986 40774 72038 40826
rect 72050 40774 72102 40826
rect 72114 40774 72166 40826
rect 65892 40672 65944 40724
rect 66076 40672 66128 40724
rect 66352 40672 66404 40724
rect 69480 40604 69532 40656
rect 65524 40536 65576 40588
rect 66076 40536 66128 40588
rect 70032 40468 70084 40520
rect 74210 40230 74262 40282
rect 74274 40230 74326 40282
rect 74338 40230 74390 40282
rect 74402 40230 74454 40282
rect 74466 40230 74518 40282
rect 65064 40128 65116 40180
rect 66352 40128 66404 40180
rect 64696 39992 64748 40044
rect 65524 39992 65576 40044
rect 71858 39686 71910 39738
rect 71922 39686 71974 39738
rect 71986 39686 72038 39738
rect 72050 39686 72102 39738
rect 72114 39686 72166 39738
rect 66168 39584 66220 39636
rect 63500 39516 63552 39568
rect 68376 39380 68428 39432
rect 74210 39142 74262 39194
rect 74274 39142 74326 39194
rect 74338 39142 74390 39194
rect 74402 39142 74454 39194
rect 74466 39142 74518 39194
rect 64052 38700 64104 38752
rect 63868 38632 63920 38684
rect 71858 38598 71910 38650
rect 71922 38598 71974 38650
rect 71986 38598 72038 38650
rect 72050 38598 72102 38650
rect 72114 38598 72166 38650
rect 65708 38539 65760 38548
rect 65708 38505 65717 38539
rect 65717 38505 65751 38539
rect 65751 38505 65760 38539
rect 65708 38496 65760 38505
rect 68192 38292 68244 38344
rect 74210 38054 74262 38106
rect 74274 38054 74326 38106
rect 74338 38054 74390 38106
rect 74402 38054 74454 38106
rect 74466 38054 74518 38106
rect 63500 37952 63552 38004
rect 65616 37952 65668 38004
rect 63500 37816 63552 37868
rect 63684 37816 63736 37868
rect 66904 37748 66956 37800
rect 71858 37510 71910 37562
rect 71922 37510 71974 37562
rect 71986 37510 72038 37562
rect 72050 37510 72102 37562
rect 72114 37510 72166 37562
rect 63684 37340 63736 37392
rect 74210 36966 74262 37018
rect 74274 36966 74326 37018
rect 74338 36966 74390 37018
rect 74402 36966 74454 37018
rect 74466 36966 74518 37018
rect 64512 36524 64564 36576
rect 71858 36422 71910 36474
rect 71922 36422 71974 36474
rect 71986 36422 72038 36474
rect 72050 36422 72102 36474
rect 72114 36422 72166 36474
rect 65524 36320 65576 36372
rect 65432 36116 65484 36168
rect 65524 36116 65576 36168
rect 66076 36116 66128 36168
rect 68284 36116 68336 36168
rect 74210 35878 74262 35930
rect 74274 35878 74326 35930
rect 74338 35878 74390 35930
rect 74402 35878 74454 35930
rect 74466 35878 74518 35930
rect 66996 35819 67048 35828
rect 66996 35785 67005 35819
rect 67005 35785 67039 35819
rect 67039 35785 67048 35819
rect 66996 35776 67048 35785
rect 65708 35683 65760 35692
rect 65708 35649 65717 35683
rect 65717 35649 65751 35683
rect 65751 35649 65760 35683
rect 65708 35640 65760 35649
rect 71858 35334 71910 35386
rect 71922 35334 71974 35386
rect 71986 35334 72038 35386
rect 72050 35334 72102 35386
rect 72114 35334 72166 35386
rect 63684 35164 63736 35216
rect 65432 35164 65484 35216
rect 66628 35139 66680 35148
rect 66628 35105 66637 35139
rect 66637 35105 66671 35139
rect 66671 35105 66680 35139
rect 66628 35096 66680 35105
rect 65432 35028 65484 35080
rect 74210 34790 74262 34842
rect 74274 34790 74326 34842
rect 74338 34790 74390 34842
rect 74402 34790 74454 34842
rect 74466 34790 74518 34842
rect 65340 34688 65392 34740
rect 65340 34552 65392 34604
rect 67916 34552 67968 34604
rect 67364 34484 67416 34536
rect 71858 34246 71910 34298
rect 71922 34246 71974 34298
rect 71986 34246 72038 34298
rect 72050 34246 72102 34298
rect 72114 34246 72166 34298
rect 65248 34144 65300 34196
rect 64696 33940 64748 33992
rect 67456 33940 67508 33992
rect 74210 33702 74262 33754
rect 74274 33702 74326 33754
rect 74338 33702 74390 33754
rect 74402 33702 74454 33754
rect 74466 33702 74518 33754
rect 63684 33124 63736 33176
rect 71858 33158 71910 33210
rect 71922 33158 71974 33210
rect 71986 33158 72038 33210
rect 72050 33158 72102 33210
rect 72114 33158 72166 33210
rect 65156 33056 65208 33108
rect 66628 32852 66680 32904
rect 74210 32614 74262 32666
rect 74274 32614 74326 32666
rect 74338 32614 74390 32666
rect 74402 32614 74454 32666
rect 74466 32614 74518 32666
rect 69572 32376 69624 32428
rect 71858 32070 71910 32122
rect 71922 32070 71974 32122
rect 71986 32070 72038 32122
rect 72050 32070 72102 32122
rect 72114 32070 72166 32122
rect 64972 31968 65024 32020
rect 64236 31696 64288 31748
rect 63684 31560 63736 31612
rect 64512 31696 64564 31748
rect 64604 31714 64656 31766
rect 66812 31764 66864 31816
rect 64236 31492 64288 31544
rect 64420 31492 64472 31544
rect 64512 31492 64564 31544
rect 63684 31424 63736 31476
rect 74210 31526 74262 31578
rect 74274 31526 74326 31578
rect 74338 31526 74390 31578
rect 74402 31526 74454 31578
rect 74466 31526 74518 31578
rect 71858 30982 71910 31034
rect 71922 30982 71974 31034
rect 71986 30982 72038 31034
rect 72050 30982 72102 31034
rect 72114 30982 72166 31034
rect 65064 30880 65116 30932
rect 65156 30812 65208 30864
rect 66720 30676 66772 30728
rect 74210 30438 74262 30490
rect 74274 30438 74326 30490
rect 74338 30438 74390 30490
rect 74402 30438 74454 30490
rect 74466 30438 74518 30490
rect 64420 30336 64472 30388
rect 64972 30336 65024 30388
rect 68008 30132 68060 30184
rect 71858 29894 71910 29946
rect 71922 29894 71974 29946
rect 71986 29894 72038 29946
rect 72050 29894 72102 29946
rect 72114 29894 72166 29946
rect 66168 29792 66220 29844
rect 68468 29724 68520 29776
rect 66352 29631 66404 29640
rect 66352 29597 66361 29631
rect 66361 29597 66395 29631
rect 66395 29597 66404 29631
rect 66352 29588 66404 29597
rect 74210 29350 74262 29402
rect 74274 29350 74326 29402
rect 74338 29350 74390 29402
rect 74402 29350 74454 29402
rect 74466 29350 74518 29402
rect 71858 28806 71910 28858
rect 71922 28806 71974 28858
rect 71986 28806 72038 28858
rect 72050 28806 72102 28858
rect 72114 28806 72166 28858
rect 65156 28636 65208 28688
rect 65708 28475 65760 28484
rect 65708 28441 65717 28475
rect 65717 28441 65751 28475
rect 65751 28441 65760 28475
rect 65708 28432 65760 28441
rect 65524 28364 65576 28416
rect 74210 28262 74262 28314
rect 74274 28262 74326 28314
rect 74338 28262 74390 28314
rect 74402 28262 74454 28314
rect 74466 28262 74518 28314
rect 65340 28160 65392 28212
rect 66260 27999 66312 28008
rect 66260 27965 66269 27999
rect 66269 27965 66303 27999
rect 66303 27965 66312 27999
rect 66260 27956 66312 27965
rect 64420 27888 64472 27940
rect 70124 27820 70176 27872
rect 71858 27718 71910 27770
rect 71922 27718 71974 27770
rect 71986 27718 72038 27770
rect 72050 27718 72102 27770
rect 72114 27718 72166 27770
rect 65432 27548 65484 27600
rect 67272 27412 67324 27464
rect 74210 27174 74262 27226
rect 74274 27174 74326 27226
rect 74338 27174 74390 27226
rect 74402 27174 74454 27226
rect 74466 27174 74518 27226
rect 66536 27004 66588 27056
rect 65616 26936 65668 26988
rect 65156 26732 65208 26784
rect 66628 26732 66680 26784
rect 66812 26732 66864 26784
rect 71858 26630 71910 26682
rect 71922 26630 71974 26682
rect 71986 26630 72038 26682
rect 72050 26630 72102 26682
rect 72114 26630 72166 26682
rect 64880 26528 64932 26580
rect 66720 26324 66772 26376
rect 74210 26086 74262 26138
rect 74274 26086 74326 26138
rect 74338 26086 74390 26138
rect 74402 26086 74454 26138
rect 74466 26086 74518 26138
rect 69940 25644 69992 25696
rect 71858 25542 71910 25594
rect 71922 25542 71974 25594
rect 71986 25542 72038 25594
rect 72050 25542 72102 25594
rect 72114 25542 72166 25594
rect 64604 25440 64656 25492
rect 64604 25236 64656 25288
rect 65432 25236 65484 25288
rect 74210 24998 74262 25050
rect 74274 24998 74326 25050
rect 74338 24998 74390 25050
rect 74402 24998 74454 25050
rect 74466 24998 74518 25050
rect 66076 24803 66128 24812
rect 66076 24769 66085 24803
rect 66085 24769 66119 24803
rect 66119 24769 66128 24803
rect 66076 24760 66128 24769
rect 66168 24692 66220 24744
rect 65432 24556 65484 24608
rect 66076 24556 66128 24608
rect 71858 24454 71910 24506
rect 71922 24454 71974 24506
rect 71986 24454 72038 24506
rect 72050 24454 72102 24506
rect 72114 24454 72166 24506
rect 65892 24395 65944 24404
rect 65892 24361 65901 24395
rect 65901 24361 65935 24395
rect 65935 24361 65944 24395
rect 65892 24352 65944 24361
rect 65984 24352 66036 24404
rect 64880 24284 64932 24336
rect 67272 24284 67324 24336
rect 67640 24284 67692 24336
rect 66076 24148 66128 24200
rect 67272 24191 67324 24200
rect 67272 24157 67281 24191
rect 67281 24157 67315 24191
rect 67315 24157 67324 24191
rect 67272 24148 67324 24157
rect 65892 24012 65944 24064
rect 66168 24012 66220 24064
rect 74210 23910 74262 23962
rect 74274 23910 74326 23962
rect 74338 23910 74390 23962
rect 74402 23910 74454 23962
rect 74466 23910 74518 23962
rect 65800 23808 65852 23860
rect 66444 23851 66496 23860
rect 66444 23817 66453 23851
rect 66453 23817 66487 23851
rect 66487 23817 66496 23851
rect 66444 23808 66496 23817
rect 67180 23851 67232 23860
rect 67180 23817 67189 23851
rect 67189 23817 67223 23851
rect 67223 23817 67232 23851
rect 67180 23808 67232 23817
rect 65248 23740 65300 23792
rect 66168 23740 66220 23792
rect 65340 23604 65392 23656
rect 67180 23604 67232 23656
rect 67732 23647 67784 23656
rect 67732 23613 67741 23647
rect 67741 23613 67775 23647
rect 67775 23613 67784 23647
rect 67732 23604 67784 23613
rect 67824 23536 67876 23588
rect 71858 23366 71910 23418
rect 71922 23366 71974 23418
rect 71986 23366 72038 23418
rect 72050 23366 72102 23418
rect 72114 23366 72166 23418
rect 63684 23264 63736 23316
rect 67548 23264 67600 23316
rect 66260 23196 66312 23248
rect 67272 23196 67324 23248
rect 63684 23060 63736 23112
rect 66536 23103 66588 23112
rect 66536 23069 66545 23103
rect 66545 23069 66579 23103
rect 66579 23069 66588 23103
rect 66536 23060 66588 23069
rect 67180 23103 67232 23112
rect 67180 23069 67189 23103
rect 67189 23069 67223 23103
rect 67223 23069 67232 23103
rect 67180 23060 67232 23069
rect 67640 23060 67692 23112
rect 67824 23060 67876 23112
rect 65340 22924 65392 22976
rect 74210 22822 74262 22874
rect 74274 22822 74326 22874
rect 74338 22822 74390 22874
rect 74402 22822 74454 22874
rect 74466 22822 74518 22874
rect 63500 22720 63552 22772
rect 63500 22516 63552 22568
rect 64880 22516 64932 22568
rect 66260 22559 66312 22568
rect 66260 22525 66269 22559
rect 66269 22525 66303 22559
rect 66303 22525 66312 22559
rect 66260 22516 66312 22525
rect 64512 22312 64564 22364
rect 64604 22312 64656 22364
rect 64880 22312 64932 22364
rect 71858 22278 71910 22330
rect 71922 22278 71974 22330
rect 71986 22278 72038 22330
rect 72050 22278 72102 22330
rect 72114 22278 72166 22330
rect 64420 22108 64472 22160
rect 64512 22108 64564 22160
rect 64604 22040 64656 22092
rect 64420 21972 64472 22024
rect 64880 21972 64932 22024
rect 74210 21734 74262 21786
rect 74274 21734 74326 21786
rect 74338 21734 74390 21786
rect 74402 21734 74454 21786
rect 74466 21734 74518 21786
rect 70216 21360 70268 21412
rect 63500 21292 63552 21344
rect 63500 21192 63552 21244
rect 71858 21190 71910 21242
rect 71922 21190 71974 21242
rect 71986 21190 72038 21242
rect 72050 21190 72102 21242
rect 72114 21190 72166 21242
rect 74210 20646 74262 20698
rect 74274 20646 74326 20698
rect 74338 20646 74390 20698
rect 74402 20646 74454 20698
rect 74466 20646 74518 20698
rect 71858 20102 71910 20154
rect 71922 20102 71974 20154
rect 71986 20102 72038 20154
rect 72050 20102 72102 20154
rect 72114 20102 72166 20154
rect 74210 19558 74262 19610
rect 74274 19558 74326 19610
rect 74338 19558 74390 19610
rect 74402 19558 74454 19610
rect 74466 19558 74518 19610
rect 64880 19252 64932 19304
rect 66260 19116 66312 19168
rect 71858 19014 71910 19066
rect 71922 19014 71974 19066
rect 71986 19014 72038 19066
rect 72050 19014 72102 19066
rect 72114 19014 72166 19066
rect 67824 18912 67876 18964
rect 74210 18470 74262 18522
rect 74274 18470 74326 18522
rect 74338 18470 74390 18522
rect 74402 18470 74454 18522
rect 74466 18470 74518 18522
rect 63684 18028 63736 18080
rect 64880 18028 64932 18080
rect 71858 17926 71910 17978
rect 71922 17926 71974 17978
rect 71986 17926 72038 17978
rect 72050 17926 72102 17978
rect 72114 17926 72166 17978
rect 64604 17552 64656 17604
rect 65064 17552 65116 17604
rect 64144 17416 64196 17468
rect 64604 17416 64656 17468
rect 74210 17382 74262 17434
rect 74274 17382 74326 17434
rect 74338 17382 74390 17434
rect 74402 17382 74454 17434
rect 74466 17382 74518 17434
rect 66536 17212 66588 17264
rect 66812 17212 66864 17264
rect 71858 16838 71910 16890
rect 71922 16838 71974 16890
rect 71986 16838 72038 16890
rect 72050 16838 72102 16890
rect 72114 16838 72166 16890
rect 65892 16736 65944 16788
rect 65984 16600 66036 16652
rect 74210 16294 74262 16346
rect 74274 16294 74326 16346
rect 74338 16294 74390 16346
rect 74402 16294 74454 16346
rect 74466 16294 74518 16346
rect 71858 15750 71910 15802
rect 71922 15750 71974 15802
rect 71986 15750 72038 15802
rect 72050 15750 72102 15802
rect 72114 15750 72166 15802
rect 63592 15580 63644 15632
rect 74210 15206 74262 15258
rect 74274 15206 74326 15258
rect 74338 15206 74390 15258
rect 74402 15206 74454 15258
rect 74466 15206 74518 15258
rect 66812 14764 66864 14816
rect 71858 14662 71910 14714
rect 71922 14662 71974 14714
rect 71986 14662 72038 14714
rect 72050 14662 72102 14714
rect 72114 14662 72166 14714
rect 65248 14356 65300 14408
rect 74210 14118 74262 14170
rect 74274 14118 74326 14170
rect 74338 14118 74390 14170
rect 74402 14118 74454 14170
rect 74466 14118 74518 14170
rect 63592 13676 63644 13728
rect 71858 13574 71910 13626
rect 71922 13574 71974 13626
rect 71986 13574 72038 13626
rect 72050 13574 72102 13626
rect 72114 13574 72166 13626
rect 74210 13030 74262 13082
rect 74274 13030 74326 13082
rect 74338 13030 74390 13082
rect 74402 13030 74454 13082
rect 74466 13030 74518 13082
rect 66076 12588 66128 12640
rect 64880 12452 64932 12504
rect 71858 12486 71910 12538
rect 71922 12486 71974 12538
rect 71986 12486 72038 12538
rect 72050 12486 72102 12538
rect 72114 12486 72166 12538
rect 63684 12384 63736 12436
rect 65064 12384 65116 12436
rect 63960 11976 64012 12028
rect 64788 11976 64840 12028
rect 74210 11942 74262 11994
rect 74274 11942 74326 11994
rect 74338 11942 74390 11994
rect 74402 11942 74454 11994
rect 74466 11942 74518 11994
rect 64604 11840 64656 11892
rect 64788 11840 64840 11892
rect 65064 11840 65116 11892
rect 65340 11840 65392 11892
rect 63592 11500 63644 11552
rect 71858 11398 71910 11450
rect 71922 11398 71974 11450
rect 71986 11398 72038 11450
rect 72050 11398 72102 11450
rect 72114 11398 72166 11450
rect 74210 10854 74262 10906
rect 74274 10854 74326 10906
rect 74338 10854 74390 10906
rect 74402 10854 74454 10906
rect 74466 10854 74518 10906
rect 63592 10292 63644 10344
rect 66536 10684 66588 10736
rect 67180 10684 67232 10736
rect 66812 10548 66864 10600
rect 67180 10548 67232 10600
rect 71858 10310 71910 10362
rect 71922 10310 71974 10362
rect 71986 10310 72038 10362
rect 72050 10310 72102 10362
rect 72114 10310 72166 10362
rect 66812 10208 66864 10260
rect 63500 10004 63552 10056
rect 74210 9766 74262 9818
rect 74274 9766 74326 9818
rect 74338 9766 74390 9818
rect 74402 9766 74454 9818
rect 74466 9766 74518 9818
rect 71858 9222 71910 9274
rect 71922 9222 71974 9274
rect 71986 9222 72038 9274
rect 72050 9222 72102 9274
rect 72114 9222 72166 9274
rect 65432 9120 65484 9172
rect 65432 8984 65484 9036
rect 65984 8984 66036 9036
rect 66076 8780 66128 8832
rect 74210 8678 74262 8730
rect 74274 8678 74326 8730
rect 74338 8678 74390 8730
rect 74402 8678 74454 8730
rect 74466 8678 74518 8730
rect 66444 8236 66496 8288
rect 71858 8134 71910 8186
rect 71922 8134 71974 8186
rect 71986 8134 72038 8186
rect 72050 8134 72102 8186
rect 72114 8134 72166 8186
rect 66444 8032 66496 8084
rect 66904 8032 66956 8084
rect 67732 8032 67784 8084
rect 50712 7828 50764 7880
rect 62488 7828 62540 7880
rect 64236 7896 64288 7948
rect 63224 7828 63276 7880
rect 67916 7896 67968 7948
rect 68652 7896 68704 7948
rect 63408 7760 63460 7812
rect 66352 7760 66404 7812
rect 66444 7760 66496 7812
rect 66536 7760 66588 7812
rect 66996 7760 67048 7812
rect 35992 7692 36044 7744
rect 64052 7692 64104 7744
rect 36084 7624 36136 7676
rect 64144 7624 64196 7676
rect 32956 7556 33008 7608
rect 63684 7556 63736 7608
rect 58992 7488 59044 7540
rect 74210 7590 74262 7642
rect 74274 7590 74326 7642
rect 74338 7590 74390 7642
rect 74402 7590 74454 7642
rect 74466 7590 74518 7642
rect 64788 7488 64840 7540
rect 69204 7531 69256 7540
rect 69204 7497 69213 7531
rect 69213 7497 69247 7531
rect 69247 7497 69256 7531
rect 69204 7488 69256 7497
rect 60004 7352 60056 7404
rect 65800 7352 65852 7404
rect 66536 7395 66588 7404
rect 66536 7361 66545 7395
rect 66545 7361 66579 7395
rect 66579 7361 66588 7395
rect 66536 7352 66588 7361
rect 67088 7352 67140 7404
rect 58900 7284 58952 7336
rect 65432 7284 65484 7336
rect 59084 7216 59136 7268
rect 65984 7216 66036 7268
rect 59544 7148 59596 7200
rect 66812 7148 66864 7200
rect 59268 7080 59320 7132
rect 65156 7080 65208 7132
rect 59728 7012 59780 7064
rect 63960 7012 64012 7064
rect 71858 7046 71910 7098
rect 71922 7046 71974 7098
rect 71986 7046 72038 7098
rect 72050 7046 72102 7098
rect 72114 7046 72166 7098
rect 59360 6944 59412 6996
rect 65340 6944 65392 6996
rect 66536 6987 66588 6996
rect 66536 6953 66545 6987
rect 66545 6953 66579 6987
rect 66579 6953 66588 6987
rect 66536 6944 66588 6953
rect 69204 6987 69256 6996
rect 69204 6953 69213 6987
rect 69213 6953 69247 6987
rect 69247 6953 69256 6987
rect 69204 6944 69256 6953
rect 61200 6876 61252 6928
rect 63500 6876 63552 6928
rect 48136 6808 48188 6860
rect 36636 6740 36688 6792
rect 64236 6740 64288 6792
rect 64604 6808 64656 6860
rect 67456 6808 67508 6860
rect 69296 6740 69348 6792
rect 35164 6672 35216 6724
rect 62856 6672 62908 6724
rect 51448 6604 51500 6656
rect 68468 6604 68520 6656
rect 33692 6536 33744 6588
rect 64512 6536 64564 6588
rect 30472 6468 30524 6520
rect 74210 6502 74262 6554
rect 74274 6502 74326 6554
rect 74338 6502 74390 6554
rect 74402 6502 74454 6554
rect 74466 6502 74518 6554
rect 30288 6400 30340 6452
rect 31024 6332 31076 6384
rect 52276 6400 52328 6452
rect 64420 6400 64472 6452
rect 65892 6400 65944 6452
rect 66536 6443 66588 6452
rect 66536 6409 66545 6443
rect 66545 6409 66579 6443
rect 66579 6409 66588 6443
rect 66536 6400 66588 6409
rect 69204 6443 69256 6452
rect 69204 6409 69213 6443
rect 69213 6409 69247 6443
rect 69247 6409 69256 6443
rect 69204 6400 69256 6409
rect 53104 6332 53156 6384
rect 62764 6332 62816 6384
rect 62856 6332 62908 6384
rect 69388 6332 69440 6384
rect 67180 6264 67232 6316
rect 53104 6196 53156 6248
rect 56600 6196 56652 6248
rect 64880 6196 64932 6248
rect 47308 6128 47360 6180
rect 65524 6128 65576 6180
rect 65892 6128 65944 6180
rect 69020 6128 69072 6180
rect 53288 6060 53340 6112
rect 61476 6060 61528 6112
rect 62764 6060 62816 6112
rect 64052 6060 64104 6112
rect 64236 6060 64288 6112
rect 69572 6060 69624 6112
rect 71858 5958 71910 6010
rect 71922 5958 71974 6010
rect 71986 5958 72038 6010
rect 72050 5958 72102 6010
rect 72114 5958 72166 6010
rect 50712 5899 50764 5908
rect 50712 5865 50721 5899
rect 50721 5865 50755 5899
rect 50755 5865 50764 5899
rect 50712 5856 50764 5865
rect 51448 5899 51500 5908
rect 51448 5865 51457 5899
rect 51457 5865 51491 5899
rect 51491 5865 51500 5899
rect 51448 5856 51500 5865
rect 52276 5856 52328 5908
rect 53288 5899 53340 5908
rect 53288 5865 53297 5899
rect 53297 5865 53331 5899
rect 53331 5865 53340 5899
rect 53288 5856 53340 5865
rect 42708 5831 42760 5840
rect 42708 5797 42717 5831
rect 42717 5797 42751 5831
rect 42751 5797 42760 5831
rect 42708 5788 42760 5797
rect 44732 5831 44784 5840
rect 44732 5797 44741 5831
rect 44741 5797 44775 5831
rect 44775 5797 44784 5831
rect 44732 5788 44784 5797
rect 59176 5899 59228 5908
rect 59176 5865 59185 5899
rect 59185 5865 59219 5899
rect 59219 5865 59228 5899
rect 59176 5856 59228 5865
rect 59728 5899 59780 5908
rect 59728 5865 59737 5899
rect 59737 5865 59771 5899
rect 59771 5865 59780 5899
rect 59728 5856 59780 5865
rect 60740 5856 60792 5908
rect 61200 5899 61252 5908
rect 61200 5865 61209 5899
rect 61209 5865 61243 5899
rect 61243 5865 61252 5899
rect 61200 5856 61252 5865
rect 61292 5856 61344 5908
rect 63500 5856 63552 5908
rect 63592 5899 63644 5908
rect 63592 5865 63601 5899
rect 63601 5865 63635 5899
rect 63635 5865 63644 5899
rect 63592 5856 63644 5865
rect 64788 5856 64840 5908
rect 66536 5899 66588 5908
rect 66536 5865 66545 5899
rect 66545 5865 66579 5899
rect 66579 5865 66588 5899
rect 66536 5856 66588 5865
rect 69204 5899 69256 5908
rect 69204 5865 69213 5899
rect 69213 5865 69247 5899
rect 69247 5865 69256 5899
rect 69204 5856 69256 5865
rect 31116 5652 31168 5704
rect 34796 5652 34848 5704
rect 35900 5652 35952 5704
rect 41512 5652 41564 5704
rect 42524 5695 42576 5704
rect 42524 5661 42533 5695
rect 42533 5661 42567 5695
rect 42567 5661 42576 5695
rect 42524 5652 42576 5661
rect 33232 5584 33284 5636
rect 45560 5652 45612 5704
rect 29828 5516 29880 5568
rect 36176 5516 36228 5568
rect 47216 5516 47268 5568
rect 49056 5652 49108 5704
rect 50804 5695 50856 5704
rect 50804 5661 50813 5695
rect 50813 5661 50847 5695
rect 50847 5661 50856 5695
rect 50804 5652 50856 5661
rect 51264 5652 51316 5704
rect 51724 5652 51776 5704
rect 52736 5652 52788 5704
rect 51172 5584 51224 5636
rect 55220 5695 55272 5704
rect 55220 5661 55229 5695
rect 55229 5661 55263 5695
rect 55263 5661 55272 5695
rect 55220 5652 55272 5661
rect 55956 5695 56008 5704
rect 55956 5661 55965 5695
rect 55965 5661 55999 5695
rect 55999 5661 56008 5695
rect 55956 5652 56008 5661
rect 56600 5695 56652 5704
rect 56600 5661 56609 5695
rect 56609 5661 56643 5695
rect 56643 5661 56652 5695
rect 56600 5652 56652 5661
rect 56692 5695 56744 5704
rect 56692 5661 56701 5695
rect 56701 5661 56735 5695
rect 56735 5661 56744 5695
rect 56692 5652 56744 5661
rect 57336 5763 57388 5772
rect 57336 5729 57345 5763
rect 57345 5729 57379 5763
rect 57379 5729 57388 5763
rect 57336 5720 57388 5729
rect 65248 5788 65300 5840
rect 65800 5788 65852 5840
rect 66168 5788 66220 5840
rect 60832 5720 60884 5772
rect 64052 5720 64104 5772
rect 70216 5720 70268 5772
rect 64696 5652 64748 5704
rect 64788 5652 64840 5704
rect 66996 5652 67048 5704
rect 62856 5584 62908 5636
rect 62304 5559 62356 5568
rect 62304 5525 62313 5559
rect 62313 5525 62347 5559
rect 62347 5525 62356 5559
rect 62304 5516 62356 5525
rect 65892 5584 65944 5636
rect 66168 5584 66220 5636
rect 67548 5584 67600 5636
rect 63500 5516 63552 5568
rect 67732 5516 67784 5568
rect 4210 5414 4262 5466
rect 4274 5414 4326 5466
rect 4338 5414 4390 5466
rect 4402 5414 4454 5466
rect 4466 5414 4518 5466
rect 14210 5414 14262 5466
rect 14274 5414 14326 5466
rect 14338 5414 14390 5466
rect 14402 5414 14454 5466
rect 14466 5414 14518 5466
rect 24210 5414 24262 5466
rect 24274 5414 24326 5466
rect 24338 5414 24390 5466
rect 24402 5414 24454 5466
rect 24466 5414 24518 5466
rect 34210 5414 34262 5466
rect 34274 5414 34326 5466
rect 34338 5414 34390 5466
rect 34402 5414 34454 5466
rect 34466 5414 34518 5466
rect 44210 5414 44262 5466
rect 44274 5414 44326 5466
rect 44338 5414 44390 5466
rect 44402 5414 44454 5466
rect 44466 5414 44518 5466
rect 54210 5414 54262 5466
rect 54274 5414 54326 5466
rect 54338 5414 54390 5466
rect 54402 5414 54454 5466
rect 54466 5414 54518 5466
rect 64210 5414 64262 5466
rect 64274 5414 64326 5466
rect 64338 5414 64390 5466
rect 64402 5414 64454 5466
rect 64466 5414 64518 5466
rect 74210 5414 74262 5466
rect 74274 5414 74326 5466
rect 74338 5414 74390 5466
rect 74402 5414 74454 5466
rect 74466 5414 74518 5466
rect 30748 5287 30800 5296
rect 30748 5253 30757 5287
rect 30757 5253 30791 5287
rect 30791 5253 30800 5287
rect 30748 5244 30800 5253
rect 31024 5355 31076 5364
rect 31024 5321 31033 5355
rect 31033 5321 31067 5355
rect 31067 5321 31076 5355
rect 31024 5312 31076 5321
rect 31392 5312 31444 5364
rect 36452 5312 36504 5364
rect 31116 5287 31168 5296
rect 31116 5253 31125 5287
rect 31125 5253 31159 5287
rect 31159 5253 31168 5287
rect 31116 5244 31168 5253
rect 31208 5244 31260 5296
rect 32404 5244 32456 5296
rect 32588 5244 32640 5296
rect 45284 5312 45336 5364
rect 45376 5312 45428 5364
rect 48504 5312 48556 5364
rect 59084 5312 59136 5364
rect 65984 5312 66036 5364
rect 66260 5312 66312 5364
rect 66536 5355 66588 5364
rect 66536 5321 66545 5355
rect 66545 5321 66579 5355
rect 66579 5321 66588 5355
rect 66536 5312 66588 5321
rect 69204 5355 69256 5364
rect 69204 5321 69213 5355
rect 69213 5321 69247 5355
rect 69247 5321 69256 5355
rect 69204 5312 69256 5321
rect 30564 5176 30616 5228
rect 30932 5176 30984 5228
rect 31300 5176 31352 5228
rect 31668 5176 31720 5228
rect 32496 5219 32548 5228
rect 32496 5185 32505 5219
rect 32505 5185 32539 5219
rect 32539 5185 32548 5219
rect 32496 5176 32548 5185
rect 34612 5176 34664 5228
rect 47216 5244 47268 5296
rect 47308 5287 47360 5296
rect 47308 5253 47317 5287
rect 47317 5253 47351 5287
rect 47351 5253 47360 5287
rect 47308 5244 47360 5253
rect 61752 5244 61804 5296
rect 62304 5244 62356 5296
rect 62396 5244 62448 5296
rect 63868 5244 63920 5296
rect 32312 5151 32364 5160
rect 32312 5117 32321 5151
rect 32321 5117 32355 5151
rect 32355 5117 32364 5151
rect 32312 5108 32364 5117
rect 32404 5108 32456 5160
rect 43904 5108 43956 5160
rect 44916 5108 44968 5160
rect 45560 5151 45612 5160
rect 45560 5117 45569 5151
rect 45569 5117 45603 5151
rect 45603 5117 45612 5151
rect 45560 5108 45612 5117
rect 65340 5176 65392 5228
rect 47584 5151 47636 5160
rect 47584 5117 47593 5151
rect 47593 5117 47627 5151
rect 47627 5117 47636 5151
rect 47584 5108 47636 5117
rect 48412 5151 48464 5160
rect 48412 5117 48421 5151
rect 48421 5117 48455 5151
rect 48455 5117 48464 5151
rect 48412 5108 48464 5117
rect 48504 5108 48556 5160
rect 52460 5108 52512 5160
rect 29920 5083 29972 5092
rect 29920 5049 29929 5083
rect 29929 5049 29963 5083
rect 29963 5049 29972 5083
rect 29920 5040 29972 5049
rect 32220 5040 32272 5092
rect 30840 4972 30892 5024
rect 31392 4972 31444 5024
rect 34704 5015 34756 5024
rect 34704 4981 34713 5015
rect 34713 4981 34747 5015
rect 34747 4981 34756 5015
rect 34704 4972 34756 4981
rect 35164 5015 35216 5024
rect 35164 4981 35173 5015
rect 35173 4981 35207 5015
rect 35207 4981 35216 5015
rect 35164 4972 35216 4981
rect 35532 4972 35584 5024
rect 36452 4972 36504 5024
rect 43904 4972 43956 5024
rect 45468 5083 45520 5092
rect 45468 5049 45477 5083
rect 45477 5049 45511 5083
rect 45511 5049 45520 5083
rect 45468 5040 45520 5049
rect 60280 5108 60332 5160
rect 62764 5108 62816 5160
rect 45744 4972 45796 5024
rect 49056 4972 49108 5024
rect 61108 5040 61160 5092
rect 63776 5040 63828 5092
rect 58900 4972 58952 5024
rect 59176 5015 59228 5024
rect 59176 4981 59185 5015
rect 59185 4981 59219 5015
rect 59219 4981 59228 5015
rect 59176 4972 59228 4981
rect 60740 4972 60792 5024
rect 63592 5015 63644 5024
rect 63592 4981 63601 5015
rect 63601 4981 63635 5015
rect 63635 4981 63644 5015
rect 63592 4972 63644 4981
rect 1858 4870 1910 4922
rect 1922 4870 1974 4922
rect 1986 4870 2038 4922
rect 2050 4870 2102 4922
rect 2114 4870 2166 4922
rect 11858 4870 11910 4922
rect 11922 4870 11974 4922
rect 11986 4870 12038 4922
rect 12050 4870 12102 4922
rect 12114 4870 12166 4922
rect 21858 4870 21910 4922
rect 21922 4870 21974 4922
rect 21986 4870 22038 4922
rect 22050 4870 22102 4922
rect 22114 4870 22166 4922
rect 31858 4870 31910 4922
rect 31922 4870 31974 4922
rect 31986 4870 32038 4922
rect 32050 4870 32102 4922
rect 32114 4870 32166 4922
rect 41858 4870 41910 4922
rect 41922 4870 41974 4922
rect 41986 4870 42038 4922
rect 42050 4870 42102 4922
rect 42114 4870 42166 4922
rect 51858 4870 51910 4922
rect 51922 4870 51974 4922
rect 51986 4870 52038 4922
rect 52050 4870 52102 4922
rect 52114 4870 52166 4922
rect 61858 4870 61910 4922
rect 61922 4870 61974 4922
rect 61986 4870 62038 4922
rect 62050 4870 62102 4922
rect 62114 4870 62166 4922
rect 71858 4870 71910 4922
rect 71922 4870 71974 4922
rect 71986 4870 72038 4922
rect 72050 4870 72102 4922
rect 72114 4870 72166 4922
rect 31208 4768 31260 4820
rect 32404 4768 32456 4820
rect 32312 4700 32364 4752
rect 29920 4632 29972 4684
rect 34060 4768 34112 4820
rect 45468 4768 45520 4820
rect 60464 4768 60516 4820
rect 62304 4768 62356 4820
rect 66536 4811 66588 4820
rect 66536 4777 66545 4811
rect 66545 4777 66579 4811
rect 66579 4777 66588 4811
rect 66536 4768 66588 4777
rect 69204 4811 69256 4820
rect 69204 4777 69213 4811
rect 69213 4777 69247 4811
rect 69247 4777 69256 4811
rect 69204 4768 69256 4777
rect 33968 4632 34020 4684
rect 34980 4632 35032 4684
rect 29368 4564 29420 4616
rect 30932 4607 30984 4616
rect 30932 4573 30941 4607
rect 30941 4573 30975 4607
rect 30975 4573 30984 4607
rect 30932 4564 30984 4573
rect 32772 4607 32824 4616
rect 32772 4573 32781 4607
rect 32781 4573 32815 4607
rect 32815 4573 32824 4607
rect 32772 4564 32824 4573
rect 32864 4564 32916 4616
rect 34612 4564 34664 4616
rect 29460 4496 29512 4548
rect 30472 4539 30524 4548
rect 30472 4505 30481 4539
rect 30481 4505 30515 4539
rect 30515 4505 30524 4539
rect 30472 4496 30524 4505
rect 30748 4539 30800 4548
rect 30748 4505 30757 4539
rect 30757 4505 30791 4539
rect 30791 4505 30800 4539
rect 30748 4496 30800 4505
rect 31116 4496 31168 4548
rect 33876 4539 33928 4548
rect 33876 4505 33885 4539
rect 33885 4505 33919 4539
rect 33919 4505 33928 4539
rect 33876 4496 33928 4505
rect 33968 4496 34020 4548
rect 35164 4564 35216 4616
rect 36268 4632 36320 4684
rect 40040 4632 40092 4684
rect 45744 4700 45796 4752
rect 46572 4632 46624 4684
rect 59268 4700 59320 4752
rect 61200 4743 61252 4752
rect 61200 4709 61209 4743
rect 61209 4709 61243 4743
rect 61243 4709 61252 4743
rect 61200 4700 61252 4709
rect 63592 4743 63644 4752
rect 63592 4709 63601 4743
rect 63601 4709 63635 4743
rect 63635 4709 63644 4743
rect 63592 4700 63644 4709
rect 63960 4700 64012 4752
rect 46940 4632 46992 4684
rect 59360 4632 59412 4684
rect 35716 4564 35768 4616
rect 36176 4564 36228 4616
rect 29828 4428 29880 4480
rect 30656 4471 30708 4480
rect 30656 4437 30665 4471
rect 30665 4437 30699 4471
rect 30699 4437 30708 4471
rect 30656 4428 30708 4437
rect 31024 4428 31076 4480
rect 31300 4471 31352 4480
rect 31300 4437 31309 4471
rect 31309 4437 31343 4471
rect 31343 4437 31352 4471
rect 31300 4428 31352 4437
rect 32956 4428 33008 4480
rect 33600 4428 33652 4480
rect 35072 4496 35124 4548
rect 44732 4564 44784 4616
rect 46848 4564 46900 4616
rect 60004 4564 60056 4616
rect 60648 4564 60700 4616
rect 53748 4496 53800 4548
rect 35164 4428 35216 4480
rect 35624 4428 35676 4480
rect 59544 4496 59596 4548
rect 60740 4496 60792 4548
rect 61476 4496 61528 4548
rect 65064 4496 65116 4548
rect 59176 4471 59228 4480
rect 59176 4437 59185 4471
rect 59185 4437 59219 4471
rect 59219 4437 59228 4471
rect 59176 4428 59228 4437
rect 59360 4428 59412 4480
rect 60832 4471 60884 4480
rect 60832 4437 60841 4471
rect 60841 4437 60875 4471
rect 60875 4437 60884 4471
rect 60832 4428 60884 4437
rect 60924 4471 60976 4480
rect 60924 4437 60933 4471
rect 60933 4437 60967 4471
rect 60967 4437 60976 4471
rect 60924 4428 60976 4437
rect 62764 4428 62816 4480
rect 70124 4428 70176 4480
rect 4210 4326 4262 4378
rect 4274 4326 4326 4378
rect 4338 4326 4390 4378
rect 4402 4326 4454 4378
rect 4466 4326 4518 4378
rect 14210 4326 14262 4378
rect 14274 4326 14326 4378
rect 14338 4326 14390 4378
rect 14402 4326 14454 4378
rect 14466 4326 14518 4378
rect 24210 4326 24262 4378
rect 24274 4326 24326 4378
rect 24338 4326 24390 4378
rect 24402 4326 24454 4378
rect 24466 4326 24518 4378
rect 34210 4326 34262 4378
rect 34274 4326 34326 4378
rect 34338 4326 34390 4378
rect 34402 4326 34454 4378
rect 34466 4326 34518 4378
rect 44210 4326 44262 4378
rect 44274 4326 44326 4378
rect 44338 4326 44390 4378
rect 44402 4326 44454 4378
rect 44466 4326 44518 4378
rect 54210 4326 54262 4378
rect 54274 4326 54326 4378
rect 54338 4326 54390 4378
rect 54402 4326 54454 4378
rect 54466 4326 54518 4378
rect 64210 4326 64262 4378
rect 64274 4326 64326 4378
rect 64338 4326 64390 4378
rect 64402 4326 64454 4378
rect 64466 4326 64518 4378
rect 74210 4326 74262 4378
rect 74274 4326 74326 4378
rect 74338 4326 74390 4378
rect 74402 4326 74454 4378
rect 74466 4326 74518 4378
rect 30656 4224 30708 4276
rect 31300 4224 31352 4276
rect 33600 4224 33652 4276
rect 34060 4224 34112 4276
rect 29368 4199 29420 4208
rect 29368 4165 29377 4199
rect 29377 4165 29411 4199
rect 29411 4165 29420 4199
rect 29368 4156 29420 4165
rect 29920 4156 29972 4208
rect 30472 4156 30524 4208
rect 32956 4199 33008 4208
rect 32956 4165 32965 4199
rect 32965 4165 32999 4199
rect 32999 4165 33008 4199
rect 32956 4156 33008 4165
rect 33968 4156 34020 4208
rect 34888 4224 34940 4276
rect 34980 4224 35032 4276
rect 35348 4267 35400 4276
rect 35348 4233 35357 4267
rect 35357 4233 35391 4267
rect 35391 4233 35400 4267
rect 35348 4224 35400 4233
rect 35808 4224 35860 4276
rect 34704 4199 34756 4208
rect 34704 4165 34713 4199
rect 34713 4165 34747 4199
rect 34747 4165 34756 4199
rect 34704 4156 34756 4165
rect 28080 4063 28132 4072
rect 28080 4029 28089 4063
rect 28089 4029 28123 4063
rect 28123 4029 28132 4063
rect 28080 4020 28132 4029
rect 29000 4020 29052 4072
rect 29828 4063 29880 4072
rect 29828 4029 29837 4063
rect 29837 4029 29871 4063
rect 29871 4029 29880 4063
rect 29828 4020 29880 4029
rect 30932 4088 30984 4140
rect 35440 4199 35492 4208
rect 35440 4165 35449 4199
rect 35449 4165 35483 4199
rect 35483 4165 35492 4199
rect 35440 4156 35492 4165
rect 35900 4156 35952 4208
rect 40776 4224 40828 4276
rect 59360 4267 59412 4276
rect 59360 4233 59369 4267
rect 59369 4233 59403 4267
rect 59403 4233 59412 4267
rect 59360 4224 59412 4233
rect 60556 4224 60608 4276
rect 60740 4224 60792 4276
rect 60832 4224 60884 4276
rect 65248 4267 65300 4276
rect 65248 4233 65257 4267
rect 65257 4233 65291 4267
rect 65291 4233 65300 4267
rect 65248 4224 65300 4233
rect 35532 4088 35584 4140
rect 35716 4131 35768 4140
rect 35716 4097 35725 4131
rect 35725 4097 35759 4131
rect 35759 4097 35768 4131
rect 35716 4088 35768 4097
rect 35808 4088 35860 4140
rect 36636 4131 36688 4140
rect 36636 4097 36645 4131
rect 36645 4097 36679 4131
rect 36679 4097 36688 4131
rect 36636 4088 36688 4097
rect 30656 4063 30708 4072
rect 30656 4029 30665 4063
rect 30665 4029 30699 4063
rect 30699 4029 30708 4063
rect 30656 4020 30708 4029
rect 31024 4020 31076 4072
rect 31668 4063 31720 4072
rect 31668 4029 31702 4063
rect 31702 4029 31720 4063
rect 31668 4020 31720 4029
rect 32312 4020 32364 4072
rect 32956 4020 33008 4072
rect 33324 4020 33376 4072
rect 33692 4020 33744 4072
rect 34060 4063 34112 4072
rect 34060 4029 34069 4063
rect 34069 4029 34103 4063
rect 34103 4029 34112 4063
rect 34060 4020 34112 4029
rect 34796 4020 34848 4072
rect 32588 3952 32640 4004
rect 36268 4063 36320 4072
rect 36268 4029 36277 4063
rect 36277 4029 36311 4063
rect 36311 4029 36320 4063
rect 36268 4020 36320 4029
rect 40224 4063 40276 4072
rect 40224 4029 40233 4063
rect 40233 4029 40267 4063
rect 40267 4029 40276 4063
rect 40224 4020 40276 4029
rect 60924 4156 60976 4208
rect 63960 4199 64012 4208
rect 63960 4165 63994 4199
rect 63994 4165 64012 4199
rect 63960 4156 64012 4165
rect 65340 4199 65392 4208
rect 65340 4165 65349 4199
rect 65349 4165 65383 4199
rect 65383 4165 65392 4199
rect 65340 4156 65392 4165
rect 40868 4088 40920 4140
rect 45376 4088 45428 4140
rect 46572 4088 46624 4140
rect 40776 4063 40828 4072
rect 40776 4029 40785 4063
rect 40785 4029 40819 4063
rect 40819 4029 40828 4063
rect 40776 4020 40828 4029
rect 27528 3927 27580 3936
rect 27528 3893 27537 3927
rect 27537 3893 27571 3927
rect 27571 3893 27580 3927
rect 27528 3884 27580 3893
rect 28632 3927 28684 3936
rect 28632 3893 28641 3927
rect 28641 3893 28675 3927
rect 28675 3893 28684 3927
rect 28632 3884 28684 3893
rect 31024 3927 31076 3936
rect 31024 3893 31033 3927
rect 31033 3893 31067 3927
rect 31067 3893 31076 3927
rect 31024 3884 31076 3893
rect 31116 3884 31168 3936
rect 31668 3884 31720 3936
rect 32220 3884 32272 3936
rect 32404 3884 32456 3936
rect 35440 3952 35492 4004
rect 35532 3952 35584 4004
rect 36452 3952 36504 4004
rect 42340 4020 42392 4072
rect 42524 4020 42576 4072
rect 40960 3952 41012 4004
rect 46296 3952 46348 4004
rect 46572 3995 46624 4004
rect 46572 3961 46581 3995
rect 46581 3961 46615 3995
rect 46615 3961 46624 3995
rect 46572 3952 46624 3961
rect 50344 4131 50396 4140
rect 50344 4097 50378 4131
rect 50378 4097 50396 4131
rect 50344 4088 50396 4097
rect 60648 4088 60700 4140
rect 65064 4088 65116 4140
rect 66536 4156 66588 4208
rect 67916 4088 67968 4140
rect 69204 4156 69256 4208
rect 48596 3952 48648 4004
rect 33140 3884 33192 3936
rect 33508 3884 33560 3936
rect 33784 3884 33836 3936
rect 34060 3884 34112 3936
rect 36176 3884 36228 3936
rect 47584 3884 47636 3936
rect 48136 3927 48188 3936
rect 48136 3893 48145 3927
rect 48145 3893 48179 3927
rect 48179 3893 48188 3927
rect 51080 3952 51132 4004
rect 51448 3952 51500 4004
rect 53380 4063 53432 4072
rect 53380 4029 53414 4063
rect 53414 4029 53432 4063
rect 53380 4020 53432 4029
rect 55036 4063 55088 4072
rect 55036 4029 55070 4063
rect 55070 4029 55088 4063
rect 55036 4020 55088 4029
rect 56508 4063 56560 4072
rect 56508 4029 56542 4063
rect 56542 4029 56560 4063
rect 56508 4020 56560 4029
rect 58256 4063 58308 4072
rect 58256 4029 58290 4063
rect 58290 4029 58308 4063
rect 58256 4020 58308 4029
rect 59176 4020 59228 4072
rect 62304 4020 62356 4072
rect 57428 3952 57480 4004
rect 61660 3952 61712 4004
rect 63868 3952 63920 4004
rect 70584 3952 70636 4004
rect 48136 3884 48188 3893
rect 52368 3884 52420 3936
rect 54024 3884 54076 3936
rect 54852 3884 54904 3936
rect 57612 3884 57664 3936
rect 58440 3927 58492 3936
rect 58440 3893 58449 3927
rect 58449 3893 58483 3927
rect 58483 3893 58492 3927
rect 58440 3884 58492 3893
rect 62672 3927 62724 3936
rect 62672 3893 62681 3927
rect 62681 3893 62715 3927
rect 62715 3893 62724 3927
rect 62672 3884 62724 3893
rect 65340 3884 65392 3936
rect 66996 3884 67048 3936
rect 69388 3884 69440 3936
rect 71412 3884 71464 3936
rect 1858 3782 1910 3834
rect 1922 3782 1974 3834
rect 1986 3782 2038 3834
rect 2050 3782 2102 3834
rect 2114 3782 2166 3834
rect 11858 3782 11910 3834
rect 11922 3782 11974 3834
rect 11986 3782 12038 3834
rect 12050 3782 12102 3834
rect 12114 3782 12166 3834
rect 21858 3782 21910 3834
rect 21922 3782 21974 3834
rect 21986 3782 22038 3834
rect 22050 3782 22102 3834
rect 22114 3782 22166 3834
rect 31858 3782 31910 3834
rect 31922 3782 31974 3834
rect 31986 3782 32038 3834
rect 32050 3782 32102 3834
rect 32114 3782 32166 3834
rect 41858 3782 41910 3834
rect 41922 3782 41974 3834
rect 41986 3782 42038 3834
rect 42050 3782 42102 3834
rect 42114 3782 42166 3834
rect 51858 3782 51910 3834
rect 51922 3782 51974 3834
rect 51986 3782 52038 3834
rect 52050 3782 52102 3834
rect 52114 3782 52166 3834
rect 61858 3782 61910 3834
rect 61922 3782 61974 3834
rect 61986 3782 62038 3834
rect 62050 3782 62102 3834
rect 62114 3782 62166 3834
rect 71858 3782 71910 3834
rect 71922 3782 71974 3834
rect 71986 3782 72038 3834
rect 72050 3782 72102 3834
rect 72114 3782 72166 3834
rect 26884 3587 26936 3596
rect 26884 3553 26893 3587
rect 26893 3553 26927 3587
rect 26927 3553 26936 3587
rect 26884 3544 26936 3553
rect 29920 3544 29972 3596
rect 30656 3544 30708 3596
rect 31693 3655 31745 3664
rect 31693 3621 31711 3655
rect 31711 3621 31745 3655
rect 31693 3612 31745 3621
rect 31392 3587 31444 3596
rect 31392 3553 31401 3587
rect 31401 3553 31435 3587
rect 31435 3553 31444 3587
rect 31392 3544 31444 3553
rect 31484 3587 31536 3596
rect 32312 3680 32364 3732
rect 33324 3680 33376 3732
rect 34796 3680 34848 3732
rect 35992 3680 36044 3732
rect 40868 3680 40920 3732
rect 41328 3680 41380 3732
rect 60648 3680 60700 3732
rect 32404 3655 32456 3664
rect 32404 3621 32413 3655
rect 32413 3621 32447 3655
rect 32447 3621 32456 3655
rect 32404 3612 32456 3621
rect 32956 3612 33008 3664
rect 33968 3612 34020 3664
rect 31484 3553 31518 3587
rect 31518 3553 31536 3587
rect 31484 3544 31536 3553
rect 27160 3519 27212 3528
rect 27160 3485 27169 3519
rect 27169 3485 27203 3519
rect 27203 3485 27212 3519
rect 27160 3476 27212 3485
rect 27988 3519 28040 3528
rect 27988 3485 27997 3519
rect 27997 3485 28031 3519
rect 28031 3485 28040 3519
rect 27988 3476 28040 3485
rect 26608 3408 26660 3460
rect 32588 3519 32640 3528
rect 29736 3451 29788 3460
rect 29736 3417 29745 3451
rect 29745 3417 29779 3451
rect 29779 3417 29788 3451
rect 29736 3408 29788 3417
rect 30288 3408 30340 3460
rect 30932 3451 30984 3460
rect 30932 3417 30941 3451
rect 30941 3417 30975 3451
rect 30975 3417 30984 3451
rect 30932 3408 30984 3417
rect 32588 3485 32597 3519
rect 32597 3485 32631 3519
rect 32631 3485 32640 3519
rect 32588 3476 32640 3485
rect 33048 3544 33100 3596
rect 33324 3519 33376 3528
rect 33324 3485 33358 3519
rect 33358 3485 33376 3519
rect 33324 3476 33376 3485
rect 33968 3476 34020 3528
rect 36084 3612 36136 3664
rect 35256 3544 35308 3596
rect 32956 3408 33008 3460
rect 27804 3383 27856 3392
rect 27804 3349 27813 3383
rect 27813 3349 27847 3383
rect 27847 3349 27856 3383
rect 27804 3340 27856 3349
rect 31392 3340 31444 3392
rect 34060 3451 34112 3460
rect 34060 3417 34094 3451
rect 34094 3417 34112 3451
rect 34060 3408 34112 3417
rect 35348 3408 35400 3460
rect 35440 3408 35492 3460
rect 40132 3544 40184 3596
rect 36360 3519 36412 3528
rect 36360 3485 36369 3519
rect 36369 3485 36403 3519
rect 36403 3485 36412 3519
rect 36360 3476 36412 3485
rect 46572 3612 46624 3664
rect 48136 3612 48188 3664
rect 51080 3612 51132 3664
rect 53104 3612 53156 3664
rect 58440 3612 58492 3664
rect 61568 3612 61620 3664
rect 45468 3476 45520 3528
rect 50988 3476 51040 3528
rect 51448 3476 51500 3528
rect 52276 3476 52328 3528
rect 57612 3519 57664 3528
rect 57612 3485 57621 3519
rect 57621 3485 57655 3519
rect 57655 3485 57664 3519
rect 57612 3476 57664 3485
rect 57796 3544 57848 3596
rect 64788 3680 64840 3732
rect 64972 3723 65024 3732
rect 64972 3689 64981 3723
rect 64981 3689 65015 3723
rect 65015 3689 65024 3723
rect 64972 3680 65024 3689
rect 66536 3723 66588 3732
rect 66536 3689 66545 3723
rect 66545 3689 66579 3723
rect 66579 3689 66588 3723
rect 66536 3680 66588 3689
rect 67916 3680 67968 3732
rect 69204 3723 69256 3732
rect 69204 3689 69213 3723
rect 69213 3689 69247 3723
rect 69247 3689 69256 3723
rect 69204 3680 69256 3689
rect 62304 3612 62356 3664
rect 63500 3612 63552 3664
rect 63960 3612 64012 3664
rect 66904 3612 66956 3664
rect 67548 3544 67600 3596
rect 61476 3476 61528 3528
rect 65432 3476 65484 3528
rect 36544 3451 36596 3460
rect 36544 3417 36553 3451
rect 36553 3417 36587 3451
rect 36587 3417 36596 3451
rect 36544 3408 36596 3417
rect 38384 3408 38436 3460
rect 33416 3340 33468 3392
rect 33600 3340 33652 3392
rect 33968 3383 34020 3392
rect 33968 3349 33977 3383
rect 33977 3349 34011 3383
rect 34011 3349 34020 3383
rect 33968 3340 34020 3349
rect 34612 3340 34664 3392
rect 34980 3383 35032 3392
rect 34980 3349 34989 3383
rect 34989 3349 35023 3383
rect 35023 3349 35032 3383
rect 34980 3340 35032 3349
rect 35072 3340 35124 3392
rect 35532 3340 35584 3392
rect 35716 3340 35768 3392
rect 40224 3408 40276 3460
rect 40316 3408 40368 3460
rect 41512 3408 41564 3460
rect 41604 3451 41656 3460
rect 41604 3417 41613 3451
rect 41613 3417 41647 3451
rect 41647 3417 41656 3451
rect 41604 3408 41656 3417
rect 42248 3408 42300 3460
rect 38844 3340 38896 3392
rect 46112 3340 46164 3392
rect 46296 3408 46348 3460
rect 48044 3408 48096 3460
rect 48136 3408 48188 3460
rect 58716 3408 58768 3460
rect 58900 3408 58952 3460
rect 52736 3340 52788 3392
rect 53012 3383 53064 3392
rect 53012 3349 53021 3383
rect 53021 3349 53055 3383
rect 53055 3349 53064 3383
rect 53012 3340 53064 3349
rect 59176 3383 59228 3392
rect 59176 3349 59185 3383
rect 59185 3349 59219 3383
rect 59219 3349 59228 3383
rect 59176 3340 59228 3349
rect 60556 3383 60608 3392
rect 60556 3349 60565 3383
rect 60565 3349 60599 3383
rect 60599 3349 60608 3383
rect 60556 3340 60608 3349
rect 60648 3340 60700 3392
rect 62580 3408 62632 3460
rect 65892 3451 65944 3460
rect 65892 3417 65901 3451
rect 65901 3417 65935 3451
rect 65935 3417 65944 3451
rect 65892 3408 65944 3417
rect 62396 3340 62448 3392
rect 69112 3340 69164 3392
rect 4210 3238 4262 3290
rect 4274 3238 4326 3290
rect 4338 3238 4390 3290
rect 4402 3238 4454 3290
rect 4466 3238 4518 3290
rect 14210 3238 14262 3290
rect 14274 3238 14326 3290
rect 14338 3238 14390 3290
rect 14402 3238 14454 3290
rect 14466 3238 14518 3290
rect 24210 3238 24262 3290
rect 24274 3238 24326 3290
rect 24338 3238 24390 3290
rect 24402 3238 24454 3290
rect 24466 3238 24518 3290
rect 34210 3238 34262 3290
rect 34274 3238 34326 3290
rect 34338 3238 34390 3290
rect 34402 3238 34454 3290
rect 34466 3238 34518 3290
rect 44210 3238 44262 3290
rect 44274 3238 44326 3290
rect 44338 3238 44390 3290
rect 44402 3238 44454 3290
rect 44466 3238 44518 3290
rect 54210 3238 54262 3290
rect 54274 3238 54326 3290
rect 54338 3238 54390 3290
rect 54402 3238 54454 3290
rect 54466 3238 54518 3290
rect 64210 3238 64262 3290
rect 64274 3238 64326 3290
rect 64338 3238 64390 3290
rect 64402 3238 64454 3290
rect 64466 3238 64518 3290
rect 74210 3238 74262 3290
rect 74274 3238 74326 3290
rect 74338 3238 74390 3290
rect 74402 3238 74454 3290
rect 74466 3238 74518 3290
rect 27988 3136 28040 3188
rect 29460 3136 29512 3188
rect 31300 3136 31352 3188
rect 32588 3136 32640 3188
rect 32772 3179 32824 3188
rect 32772 3145 32781 3179
rect 32781 3145 32815 3179
rect 32815 3145 32824 3179
rect 32772 3136 32824 3145
rect 33692 3136 33744 3188
rect 33784 3136 33836 3188
rect 39764 3136 39816 3188
rect 42248 3136 42300 3188
rect 45008 3136 45060 3188
rect 50896 3136 50948 3188
rect 50988 3136 51040 3188
rect 51724 3136 51776 3188
rect 31024 3068 31076 3120
rect 33324 3068 33376 3120
rect 34060 3068 34112 3120
rect 35532 3068 35584 3120
rect 25688 3043 25740 3052
rect 25688 3009 25697 3043
rect 25697 3009 25731 3043
rect 25731 3009 25740 3043
rect 25688 3000 25740 3009
rect 26700 3043 26752 3052
rect 26700 3009 26709 3043
rect 26709 3009 26743 3043
rect 26743 3009 26752 3043
rect 26700 3000 26752 3009
rect 28632 3000 28684 3052
rect 29920 3000 29972 3052
rect 26884 2932 26936 2984
rect 30840 3000 30892 3052
rect 31484 3000 31536 3052
rect 30104 2975 30156 2984
rect 30104 2941 30113 2975
rect 30113 2941 30147 2975
rect 30147 2941 30156 2975
rect 30104 2932 30156 2941
rect 31668 2932 31720 2984
rect 32220 2975 32272 2984
rect 32220 2941 32229 2975
rect 32229 2941 32263 2975
rect 32263 2941 32272 2975
rect 32220 2932 32272 2941
rect 30012 2864 30064 2916
rect 44916 3068 44968 3120
rect 57796 3136 57848 3188
rect 58992 3136 59044 3188
rect 59084 3179 59136 3188
rect 59084 3145 59093 3179
rect 59093 3145 59127 3179
rect 59127 3145 59136 3179
rect 59084 3136 59136 3145
rect 62488 3136 62540 3188
rect 63500 3179 63552 3188
rect 63500 3145 63509 3179
rect 63509 3145 63543 3179
rect 63543 3145 63552 3179
rect 63500 3136 63552 3145
rect 66536 3179 66588 3188
rect 66536 3145 66545 3179
rect 66545 3145 66579 3179
rect 66579 3145 66588 3179
rect 66536 3136 66588 3145
rect 69204 3179 69256 3188
rect 69204 3145 69213 3179
rect 69213 3145 69247 3179
rect 69247 3145 69256 3179
rect 69204 3136 69256 3145
rect 33140 2932 33192 2984
rect 35900 2932 35952 2984
rect 37464 2975 37516 2984
rect 37464 2941 37473 2975
rect 37473 2941 37507 2975
rect 37507 2941 37516 2975
rect 37464 2932 37516 2941
rect 37648 3043 37700 3052
rect 37648 3009 37657 3043
rect 37657 3009 37691 3043
rect 37691 3009 37700 3043
rect 37648 3000 37700 3009
rect 38200 3000 38252 3052
rect 38384 3043 38436 3052
rect 38384 3009 38393 3043
rect 38393 3009 38427 3043
rect 38427 3009 38436 3043
rect 38384 3000 38436 3009
rect 38844 3043 38896 3052
rect 38844 3009 38853 3043
rect 38853 3009 38887 3043
rect 38887 3009 38896 3043
rect 38844 3000 38896 3009
rect 39120 3043 39172 3052
rect 39120 3009 39129 3043
rect 39129 3009 39163 3043
rect 39163 3009 39172 3043
rect 39120 3000 39172 3009
rect 41328 3043 41380 3052
rect 41328 3009 41337 3043
rect 41337 3009 41371 3043
rect 41371 3009 41380 3043
rect 41328 3000 41380 3009
rect 41696 3000 41748 3052
rect 42432 3000 42484 3052
rect 37832 2975 37884 2984
rect 37832 2941 37841 2975
rect 37841 2941 37875 2975
rect 37875 2941 37884 2975
rect 37832 2932 37884 2941
rect 37924 2932 37976 2984
rect 40960 2932 41012 2984
rect 42248 2932 42300 2984
rect 29092 2796 29144 2848
rect 30564 2796 30616 2848
rect 31024 2796 31076 2848
rect 31300 2796 31352 2848
rect 33140 2796 33192 2848
rect 33416 2796 33468 2848
rect 35072 2907 35124 2916
rect 35072 2873 35081 2907
rect 35081 2873 35115 2907
rect 35115 2873 35124 2907
rect 35072 2864 35124 2873
rect 35992 2839 36044 2848
rect 35992 2805 36001 2839
rect 36001 2805 36035 2839
rect 36035 2805 36044 2839
rect 35992 2796 36044 2805
rect 36084 2796 36136 2848
rect 42524 2796 42576 2848
rect 42984 2839 43036 2848
rect 42984 2805 42993 2839
rect 42993 2805 43027 2839
rect 43027 2805 43036 2839
rect 42984 2796 43036 2805
rect 44640 3043 44692 3052
rect 44640 3009 44649 3043
rect 44649 3009 44683 3043
rect 44683 3009 44692 3043
rect 44640 3000 44692 3009
rect 45008 3000 45060 3052
rect 46112 3000 46164 3052
rect 47676 3000 47728 3052
rect 48044 3000 48096 3052
rect 59176 3068 59228 3120
rect 60556 3111 60608 3120
rect 60556 3077 60565 3111
rect 60565 3077 60599 3111
rect 60599 3077 60608 3111
rect 60556 3068 60608 3077
rect 62304 3068 62356 3120
rect 59268 3000 59320 3052
rect 59636 3043 59688 3052
rect 59636 3009 59645 3043
rect 59645 3009 59679 3043
rect 59679 3009 59688 3043
rect 59636 3000 59688 3009
rect 61568 3000 61620 3052
rect 63592 3068 63644 3120
rect 62672 3000 62724 3052
rect 69388 3043 69440 3052
rect 69388 3009 69397 3043
rect 69397 3009 69431 3043
rect 69431 3009 69440 3043
rect 69388 3000 69440 3009
rect 48136 2932 48188 2984
rect 63868 2932 63920 2984
rect 63960 2975 64012 2984
rect 63960 2941 63969 2975
rect 63969 2941 64003 2975
rect 64003 2941 64012 2975
rect 63960 2932 64012 2941
rect 64696 2932 64748 2984
rect 67640 2932 67692 2984
rect 68560 2932 68612 2984
rect 66444 2864 66496 2916
rect 45100 2796 45152 2848
rect 45468 2796 45520 2848
rect 50804 2796 50856 2848
rect 59176 2796 59228 2848
rect 62764 2796 62816 2848
rect 65524 2796 65576 2848
rect 68100 2796 68152 2848
rect 1858 2694 1910 2746
rect 1922 2694 1974 2746
rect 1986 2694 2038 2746
rect 2050 2694 2102 2746
rect 2114 2694 2166 2746
rect 11858 2694 11910 2746
rect 11922 2694 11974 2746
rect 11986 2694 12038 2746
rect 12050 2694 12102 2746
rect 12114 2694 12166 2746
rect 21858 2694 21910 2746
rect 21922 2694 21974 2746
rect 21986 2694 22038 2746
rect 22050 2694 22102 2746
rect 22114 2694 22166 2746
rect 31858 2694 31910 2746
rect 31922 2694 31974 2746
rect 31986 2694 32038 2746
rect 32050 2694 32102 2746
rect 32114 2694 32166 2746
rect 41858 2694 41910 2746
rect 41922 2694 41974 2746
rect 41986 2694 42038 2746
rect 42050 2694 42102 2746
rect 42114 2694 42166 2746
rect 51858 2694 51910 2746
rect 51922 2694 51974 2746
rect 51986 2694 52038 2746
rect 52050 2694 52102 2746
rect 52114 2694 52166 2746
rect 61858 2694 61910 2746
rect 61922 2694 61974 2746
rect 61986 2694 62038 2746
rect 62050 2694 62102 2746
rect 62114 2694 62166 2746
rect 71858 2694 71910 2746
rect 71922 2694 71974 2746
rect 71986 2694 72038 2746
rect 72050 2694 72102 2746
rect 72114 2694 72166 2746
rect 27160 2592 27212 2644
rect 30104 2592 30156 2644
rect 32220 2592 32272 2644
rect 33876 2592 33928 2644
rect 36360 2592 36412 2644
rect 37648 2592 37700 2644
rect 37832 2635 37884 2644
rect 37832 2601 37841 2635
rect 37841 2601 37875 2635
rect 37875 2601 37884 2635
rect 37832 2592 37884 2601
rect 39120 2592 39172 2644
rect 41604 2635 41656 2644
rect 41604 2601 41613 2635
rect 41613 2601 41647 2635
rect 41647 2601 41656 2635
rect 41604 2592 41656 2601
rect 41696 2635 41748 2644
rect 41696 2601 41705 2635
rect 41705 2601 41739 2635
rect 41739 2601 41748 2635
rect 41696 2592 41748 2601
rect 42432 2635 42484 2644
rect 42432 2601 42441 2635
rect 42441 2601 42475 2635
rect 42475 2601 42484 2635
rect 42432 2592 42484 2601
rect 44640 2592 44692 2644
rect 52460 2592 52512 2644
rect 48412 2524 48464 2576
rect 26240 2456 26292 2508
rect 27068 2456 27120 2508
rect 24860 2388 24912 2440
rect 27160 2388 27212 2440
rect 28172 2431 28224 2440
rect 28172 2397 28181 2431
rect 28181 2397 28215 2431
rect 28215 2397 28224 2431
rect 28172 2388 28224 2397
rect 30564 2499 30616 2508
rect 30564 2465 30573 2499
rect 30573 2465 30607 2499
rect 30607 2465 30616 2499
rect 30564 2456 30616 2465
rect 32496 2456 32548 2508
rect 33600 2456 33652 2508
rect 26792 2320 26844 2372
rect 27620 2320 27672 2372
rect 25136 2295 25188 2304
rect 25136 2261 25145 2295
rect 25145 2261 25179 2295
rect 25179 2261 25188 2295
rect 25136 2252 25188 2261
rect 25228 2252 25280 2304
rect 28448 2295 28500 2304
rect 28448 2261 28457 2295
rect 28457 2261 28491 2295
rect 28491 2261 28500 2295
rect 28448 2252 28500 2261
rect 30840 2431 30892 2440
rect 30840 2397 30849 2431
rect 30849 2397 30883 2431
rect 30883 2397 30892 2431
rect 30840 2388 30892 2397
rect 31484 2431 31536 2440
rect 31484 2397 31493 2431
rect 31493 2397 31527 2431
rect 31527 2397 31536 2431
rect 31484 2388 31536 2397
rect 33968 2388 34020 2440
rect 34980 2388 35032 2440
rect 31300 2252 31352 2304
rect 32496 2252 32548 2304
rect 35164 2252 35216 2304
rect 35992 2499 36044 2508
rect 35992 2465 36001 2499
rect 36001 2465 36035 2499
rect 36035 2465 36044 2499
rect 35992 2456 36044 2465
rect 42984 2499 43036 2508
rect 42984 2465 42993 2499
rect 42993 2465 43027 2499
rect 43027 2465 43036 2499
rect 42984 2456 43036 2465
rect 51632 2524 51684 2576
rect 37004 2388 37056 2440
rect 37740 2388 37792 2440
rect 38752 2431 38804 2440
rect 38752 2397 38761 2431
rect 38761 2397 38795 2431
rect 38795 2397 38804 2431
rect 38752 2388 38804 2397
rect 40684 2388 40736 2440
rect 41420 2388 41472 2440
rect 42708 2388 42760 2440
rect 42800 2388 42852 2440
rect 45468 2388 45520 2440
rect 46940 2388 46992 2440
rect 47400 2388 47452 2440
rect 49424 2388 49476 2440
rect 50160 2431 50212 2440
rect 50160 2397 50169 2431
rect 50169 2397 50203 2431
rect 50203 2397 50212 2431
rect 50160 2388 50212 2397
rect 56692 2456 56744 2508
rect 52644 2388 52696 2440
rect 53656 2431 53708 2440
rect 53656 2397 53665 2431
rect 53665 2397 53699 2431
rect 53699 2397 53708 2431
rect 53656 2388 53708 2397
rect 55588 2388 55640 2440
rect 56324 2431 56376 2440
rect 56324 2397 56333 2431
rect 56333 2397 56367 2431
rect 56367 2397 56376 2431
rect 56324 2388 56376 2397
rect 51632 2320 51684 2372
rect 46848 2252 46900 2304
rect 47032 2295 47084 2304
rect 47032 2261 47041 2295
rect 47041 2261 47075 2295
rect 47075 2261 47084 2295
rect 47032 2252 47084 2261
rect 48136 2295 48188 2304
rect 48136 2261 48145 2295
rect 48145 2261 48179 2295
rect 48179 2261 48188 2295
rect 48136 2252 48188 2261
rect 50804 2295 50856 2304
rect 50804 2261 50813 2295
rect 50813 2261 50847 2295
rect 50847 2261 50856 2295
rect 50804 2252 50856 2261
rect 55772 2252 55824 2304
rect 62672 2524 62724 2576
rect 63500 2635 63552 2644
rect 63500 2601 63509 2635
rect 63509 2601 63543 2635
rect 63543 2601 63552 2635
rect 63500 2592 63552 2601
rect 65892 2592 65944 2644
rect 66536 2635 66588 2644
rect 66536 2601 66545 2635
rect 66545 2601 66579 2635
rect 66579 2601 66588 2635
rect 66536 2592 66588 2601
rect 69204 2635 69256 2644
rect 69204 2601 69213 2635
rect 69213 2601 69247 2635
rect 69247 2601 69256 2635
rect 69204 2592 69256 2601
rect 63776 2524 63828 2576
rect 57520 2456 57572 2508
rect 59084 2499 59136 2508
rect 59084 2465 59093 2499
rect 59093 2465 59127 2499
rect 59127 2465 59136 2499
rect 59084 2456 59136 2465
rect 60556 2499 60608 2508
rect 60556 2465 60565 2499
rect 60565 2465 60599 2499
rect 60599 2465 60608 2499
rect 60556 2456 60608 2465
rect 61660 2456 61712 2508
rect 57428 2388 57480 2440
rect 58532 2388 58584 2440
rect 61384 2388 61436 2440
rect 62304 2431 62356 2440
rect 62304 2397 62313 2431
rect 62313 2397 62347 2431
rect 62347 2397 62356 2431
rect 62304 2388 62356 2397
rect 60096 2320 60148 2372
rect 65524 2499 65576 2508
rect 65524 2465 65533 2499
rect 65533 2465 65567 2499
rect 65567 2465 65576 2499
rect 65524 2456 65576 2465
rect 65800 2456 65852 2508
rect 68376 2499 68428 2508
rect 68376 2465 68385 2499
rect 68385 2465 68419 2499
rect 68419 2465 68428 2499
rect 68376 2456 68428 2465
rect 69848 2456 69900 2508
rect 65340 2388 65392 2440
rect 68100 2431 68152 2440
rect 68100 2397 68109 2431
rect 68109 2397 68143 2431
rect 68143 2397 68152 2431
rect 68100 2388 68152 2397
rect 69480 2431 69532 2440
rect 69480 2397 69489 2431
rect 69489 2397 69523 2431
rect 69523 2397 69532 2431
rect 69480 2388 69532 2397
rect 70676 2431 70728 2440
rect 70676 2397 70685 2431
rect 70685 2397 70719 2431
rect 70719 2397 70728 2431
rect 70676 2388 70728 2397
rect 72608 2431 72660 2440
rect 72608 2397 72617 2431
rect 72617 2397 72651 2431
rect 72651 2397 72660 2431
rect 72608 2388 72660 2397
rect 59176 2252 59228 2304
rect 60004 2252 60056 2304
rect 61016 2295 61068 2304
rect 61016 2261 61025 2295
rect 61025 2261 61059 2295
rect 61059 2261 61068 2295
rect 61016 2252 61068 2261
rect 61660 2252 61712 2304
rect 69664 2320 69716 2372
rect 62396 2252 62448 2304
rect 62580 2252 62632 2304
rect 63132 2252 63184 2304
rect 64604 2252 64656 2304
rect 70860 2252 70912 2304
rect 4210 2150 4262 2202
rect 4274 2150 4326 2202
rect 4338 2150 4390 2202
rect 4402 2150 4454 2202
rect 4466 2150 4518 2202
rect 14210 2150 14262 2202
rect 14274 2150 14326 2202
rect 14338 2150 14390 2202
rect 14402 2150 14454 2202
rect 14466 2150 14518 2202
rect 24210 2150 24262 2202
rect 24274 2150 24326 2202
rect 24338 2150 24390 2202
rect 24402 2150 24454 2202
rect 24466 2150 24518 2202
rect 34210 2150 34262 2202
rect 34274 2150 34326 2202
rect 34338 2150 34390 2202
rect 34402 2150 34454 2202
rect 34466 2150 34518 2202
rect 44210 2150 44262 2202
rect 44274 2150 44326 2202
rect 44338 2150 44390 2202
rect 44402 2150 44454 2202
rect 44466 2150 44518 2202
rect 54210 2150 54262 2202
rect 54274 2150 54326 2202
rect 54338 2150 54390 2202
rect 54402 2150 54454 2202
rect 54466 2150 54518 2202
rect 64210 2150 64262 2202
rect 64274 2150 64326 2202
rect 64338 2150 64390 2202
rect 64402 2150 64454 2202
rect 64466 2150 64518 2202
rect 74210 2150 74262 2202
rect 74274 2150 74326 2202
rect 74338 2150 74390 2202
rect 74402 2150 74454 2202
rect 74466 2150 74518 2202
rect 25688 2048 25740 2100
rect 26608 2048 26660 2100
rect 26700 2091 26752 2100
rect 26700 2057 26709 2091
rect 26709 2057 26743 2091
rect 26743 2057 26752 2091
rect 26700 2048 26752 2057
rect 27068 2091 27120 2100
rect 27068 2057 27077 2091
rect 27077 2057 27111 2091
rect 27111 2057 27120 2091
rect 27068 2048 27120 2057
rect 28448 2048 28500 2100
rect 34060 2048 34112 2100
rect 36544 2048 36596 2100
rect 37004 2091 37056 2100
rect 37004 2057 37013 2091
rect 37013 2057 37047 2091
rect 37047 2057 37056 2091
rect 37004 2048 37056 2057
rect 40684 2091 40736 2100
rect 40684 2057 40693 2091
rect 40693 2057 40727 2091
rect 40727 2057 40736 2091
rect 40684 2048 40736 2057
rect 41420 2091 41472 2100
rect 41420 2057 41429 2091
rect 41429 2057 41463 2091
rect 41463 2057 41472 2091
rect 41420 2048 41472 2057
rect 41696 2048 41748 2100
rect 44732 2048 44784 2100
rect 45100 2048 45152 2100
rect 46940 2091 46992 2100
rect 46940 2057 46949 2091
rect 46949 2057 46983 2091
rect 46983 2057 46992 2091
rect 46940 2048 46992 2057
rect 47584 2091 47636 2100
rect 47584 2057 47593 2091
rect 47593 2057 47627 2091
rect 47627 2057 47636 2091
rect 47584 2048 47636 2057
rect 49424 2091 49476 2100
rect 49424 2057 49433 2091
rect 49433 2057 49467 2091
rect 49467 2057 49476 2091
rect 49424 2048 49476 2057
rect 24676 1912 24728 1964
rect 25320 1912 25372 1964
rect 27804 1912 27856 1964
rect 29092 1955 29144 1964
rect 29092 1921 29101 1955
rect 29101 1921 29135 1955
rect 29135 1921 29144 1955
rect 29092 1912 29144 1921
rect 33968 1980 34020 2032
rect 34888 1980 34940 2032
rect 41144 1980 41196 2032
rect 48780 1980 48832 2032
rect 52644 2091 52696 2100
rect 52644 2057 52653 2091
rect 52653 2057 52687 2091
rect 52687 2057 52696 2091
rect 52644 2048 52696 2057
rect 55588 2091 55640 2100
rect 55588 2057 55597 2091
rect 55597 2057 55631 2091
rect 55631 2057 55640 2091
rect 55588 2048 55640 2057
rect 59084 2091 59136 2100
rect 59084 2057 59093 2091
rect 59093 2057 59127 2091
rect 59127 2057 59136 2091
rect 59084 2048 59136 2057
rect 59636 2048 59688 2100
rect 60556 2091 60608 2100
rect 60556 2057 60565 2091
rect 60565 2057 60599 2091
rect 60599 2057 60608 2091
rect 60556 2048 60608 2057
rect 61384 2091 61436 2100
rect 61384 2057 61393 2091
rect 61393 2057 61427 2091
rect 61427 2057 61436 2091
rect 61384 2048 61436 2057
rect 66352 2048 66404 2100
rect 66536 2091 66588 2100
rect 66536 2057 66545 2091
rect 66545 2057 66579 2091
rect 66579 2057 66588 2091
rect 66536 2048 66588 2057
rect 66996 2048 67048 2100
rect 31116 1912 31168 1964
rect 33048 1912 33100 1964
rect 33508 1955 33560 1964
rect 33508 1921 33517 1955
rect 33517 1921 33551 1955
rect 33551 1921 33560 1955
rect 33508 1912 33560 1921
rect 33876 1912 33928 1964
rect 34612 1912 34664 1964
rect 25228 1844 25280 1896
rect 25412 1887 25464 1896
rect 25412 1853 25421 1887
rect 25421 1853 25455 1887
rect 25455 1853 25464 1887
rect 25412 1844 25464 1853
rect 27528 1844 27580 1896
rect 30380 1844 30432 1896
rect 32220 1844 32272 1896
rect 34060 1844 34112 1896
rect 35624 1887 35676 1896
rect 35624 1853 35633 1887
rect 35633 1853 35667 1887
rect 35667 1853 35676 1887
rect 35624 1844 35676 1853
rect 37280 1844 37332 1896
rect 28172 1708 28224 1760
rect 30564 1708 30616 1760
rect 32496 1708 32548 1760
rect 35808 1708 35860 1760
rect 36820 1776 36872 1828
rect 39120 1844 39172 1896
rect 41236 1955 41288 1964
rect 41236 1921 41245 1955
rect 41245 1921 41279 1955
rect 41279 1921 41288 1955
rect 41236 1912 41288 1921
rect 41420 1912 41472 1964
rect 40040 1844 40092 1896
rect 42524 1912 42576 1964
rect 47032 1955 47084 1964
rect 47032 1921 47041 1955
rect 47041 1921 47075 1955
rect 47075 1921 47084 1955
rect 47032 1912 47084 1921
rect 47768 1955 47820 1964
rect 47768 1921 47777 1955
rect 47777 1921 47811 1955
rect 47811 1921 47820 1955
rect 47768 1912 47820 1921
rect 47952 1955 48004 1964
rect 47952 1921 47961 1955
rect 47961 1921 47995 1955
rect 47995 1921 48004 1955
rect 47952 1912 48004 1921
rect 50528 1955 50580 1964
rect 50528 1921 50537 1955
rect 50537 1921 50571 1955
rect 50571 1921 50580 1955
rect 50528 1912 50580 1921
rect 62396 1980 62448 2032
rect 62580 2023 62632 2032
rect 62580 1989 62589 2023
rect 62589 1989 62623 2023
rect 62623 1989 62632 2023
rect 62580 1980 62632 1989
rect 62672 1980 62724 2032
rect 65984 1980 66036 2032
rect 68008 1980 68060 2032
rect 53104 1912 53156 1964
rect 54024 1912 54076 1964
rect 41696 1708 41748 1760
rect 42432 1776 42484 1828
rect 43720 1844 43772 1896
rect 43260 1776 43312 1828
rect 46020 1844 46072 1896
rect 47860 1844 47912 1896
rect 48780 1844 48832 1896
rect 50620 1844 50672 1896
rect 51540 1844 51592 1896
rect 53380 1844 53432 1896
rect 54576 1844 54628 1896
rect 55772 1955 55824 1964
rect 55772 1921 55781 1955
rect 55781 1921 55815 1955
rect 55815 1921 55824 1955
rect 55772 1912 55824 1921
rect 57060 1912 57112 1964
rect 60004 1955 60056 1964
rect 60004 1921 60013 1955
rect 60013 1921 60047 1955
rect 60047 1921 60056 1955
rect 60004 1912 60056 1921
rect 60096 1912 60148 1964
rect 62948 1912 63000 1964
rect 56140 1844 56192 1896
rect 59820 1844 59872 1896
rect 61016 1844 61068 1896
rect 63132 1912 63184 1964
rect 63500 1955 63552 1964
rect 63500 1921 63509 1955
rect 63509 1921 63543 1955
rect 63543 1921 63552 1955
rect 63500 1912 63552 1921
rect 63684 1955 63736 1964
rect 63684 1921 63693 1955
rect 63693 1921 63727 1955
rect 63727 1921 63736 1955
rect 63684 1912 63736 1921
rect 70676 2048 70728 2100
rect 69204 2023 69256 2032
rect 69204 1989 69213 2023
rect 69213 1989 69247 2023
rect 69247 1989 69256 2023
rect 69204 1980 69256 1989
rect 70032 1980 70084 2032
rect 63224 1844 63276 1896
rect 65340 1844 65392 1896
rect 67180 1844 67232 1896
rect 70860 1955 70912 1964
rect 70860 1921 70869 1955
rect 70869 1921 70903 1955
rect 70903 1921 70912 1955
rect 70860 1912 70912 1921
rect 71412 1955 71464 1964
rect 71412 1921 71421 1955
rect 71421 1921 71455 1955
rect 71455 1921 71464 1955
rect 71412 1912 71464 1921
rect 55220 1776 55272 1828
rect 51264 1708 51316 1760
rect 58440 1751 58492 1760
rect 58440 1717 58449 1751
rect 58449 1717 58483 1751
rect 58483 1717 58492 1751
rect 58440 1708 58492 1717
rect 63408 1708 63460 1760
rect 63776 1776 63828 1828
rect 66168 1776 66220 1828
rect 71320 1844 71372 1896
rect 69388 1776 69440 1828
rect 67364 1708 67416 1760
rect 1858 1606 1910 1658
rect 1922 1606 1974 1658
rect 1986 1606 2038 1658
rect 2050 1606 2102 1658
rect 2114 1606 2166 1658
rect 11858 1606 11910 1658
rect 11922 1606 11974 1658
rect 11986 1606 12038 1658
rect 12050 1606 12102 1658
rect 12114 1606 12166 1658
rect 21858 1606 21910 1658
rect 21922 1606 21974 1658
rect 21986 1606 22038 1658
rect 22050 1606 22102 1658
rect 22114 1606 22166 1658
rect 31858 1606 31910 1658
rect 31922 1606 31974 1658
rect 31986 1606 32038 1658
rect 32050 1606 32102 1658
rect 32114 1606 32166 1658
rect 41858 1606 41910 1658
rect 41922 1606 41974 1658
rect 41986 1606 42038 1658
rect 42050 1606 42102 1658
rect 42114 1606 42166 1658
rect 51858 1606 51910 1658
rect 51922 1606 51974 1658
rect 51986 1606 52038 1658
rect 52050 1606 52102 1658
rect 52114 1606 52166 1658
rect 61858 1606 61910 1658
rect 61922 1606 61974 1658
rect 61986 1606 62038 1658
rect 62050 1606 62102 1658
rect 62114 1606 62166 1658
rect 71858 1606 71910 1658
rect 71922 1606 71974 1658
rect 71986 1606 72038 1658
rect 72050 1606 72102 1658
rect 72114 1606 72166 1658
rect 25412 1504 25464 1556
rect 29460 1504 29512 1556
rect 31484 1504 31536 1556
rect 25136 1436 25188 1488
rect 30472 1436 30524 1488
rect 32864 1504 32916 1556
rect 35624 1504 35676 1556
rect 38752 1504 38804 1556
rect 41236 1547 41288 1556
rect 41236 1513 41245 1547
rect 41245 1513 41279 1547
rect 41279 1513 41288 1547
rect 41236 1504 41288 1513
rect 59084 1547 59136 1556
rect 59084 1513 59093 1547
rect 59093 1513 59127 1547
rect 59127 1513 59136 1547
rect 59084 1504 59136 1513
rect 59176 1504 59228 1556
rect 23940 1368 23992 1420
rect 32680 1436 32732 1488
rect 34888 1436 34940 1488
rect 47584 1436 47636 1488
rect 55956 1436 56008 1488
rect 60556 1479 60608 1488
rect 60556 1445 60565 1479
rect 60565 1445 60599 1479
rect 60599 1445 60608 1479
rect 60556 1436 60608 1445
rect 62396 1436 62448 1488
rect 63500 1479 63552 1488
rect 63500 1445 63509 1479
rect 63509 1445 63543 1479
rect 63543 1445 63552 1479
rect 63500 1436 63552 1445
rect 66536 1547 66588 1556
rect 66536 1513 66545 1547
rect 66545 1513 66579 1547
rect 66579 1513 66588 1547
rect 66536 1504 66588 1513
rect 68284 1547 68336 1556
rect 68284 1513 68293 1547
rect 68293 1513 68327 1547
rect 68327 1513 68336 1547
rect 68284 1504 68336 1513
rect 69204 1547 69256 1556
rect 69204 1513 69213 1547
rect 69213 1513 69247 1547
rect 69247 1513 69256 1547
rect 69204 1504 69256 1513
rect 69480 1504 69532 1556
rect 67272 1436 67324 1488
rect 23480 1300 23532 1352
rect 25688 1343 25740 1352
rect 25688 1309 25697 1343
rect 25697 1309 25731 1343
rect 25731 1309 25740 1343
rect 25688 1300 25740 1309
rect 26884 1300 26936 1352
rect 27252 1343 27304 1352
rect 27252 1309 27261 1343
rect 27261 1309 27295 1343
rect 27295 1309 27304 1343
rect 27252 1300 27304 1309
rect 30840 1368 30892 1420
rect 33140 1368 33192 1420
rect 29828 1343 29880 1352
rect 29828 1309 29837 1343
rect 29837 1309 29871 1343
rect 29871 1309 29880 1343
rect 29828 1300 29880 1309
rect 30012 1300 30064 1352
rect 28264 1232 28316 1284
rect 28540 1232 28592 1284
rect 33968 1343 34020 1352
rect 33968 1309 33977 1343
rect 33977 1309 34011 1343
rect 34011 1309 34020 1343
rect 33968 1300 34020 1309
rect 35440 1300 35492 1352
rect 36360 1300 36412 1352
rect 38200 1343 38252 1352
rect 38200 1309 38209 1343
rect 38209 1309 38243 1343
rect 38243 1309 38252 1343
rect 38200 1300 38252 1309
rect 40500 1368 40552 1420
rect 41420 1368 41472 1420
rect 38660 1300 38712 1352
rect 39764 1343 39816 1352
rect 39764 1309 39773 1343
rect 39773 1309 39807 1343
rect 39807 1309 39816 1343
rect 39764 1300 39816 1309
rect 40040 1300 40092 1352
rect 42340 1343 42392 1352
rect 42340 1309 42349 1343
rect 42349 1309 42383 1343
rect 42383 1309 42392 1343
rect 42340 1300 42392 1309
rect 42708 1300 42760 1352
rect 43904 1300 43956 1352
rect 45192 1343 45244 1352
rect 45192 1309 45201 1343
rect 45201 1309 45235 1343
rect 45235 1309 45244 1343
rect 45192 1300 45244 1309
rect 45468 1300 45520 1352
rect 49240 1368 49292 1420
rect 58440 1368 58492 1420
rect 27620 1164 27672 1216
rect 35624 1232 35676 1284
rect 38292 1232 38344 1284
rect 39580 1232 39632 1284
rect 40960 1232 41012 1284
rect 45100 1232 45152 1284
rect 44088 1164 44140 1216
rect 44640 1164 44692 1216
rect 47492 1343 47544 1352
rect 47492 1309 47501 1343
rect 47501 1309 47535 1343
rect 47535 1309 47544 1343
rect 47492 1300 47544 1309
rect 47768 1300 47820 1352
rect 46480 1232 46532 1284
rect 48136 1164 48188 1216
rect 49608 1300 49660 1352
rect 50804 1300 50856 1352
rect 52276 1300 52328 1352
rect 53656 1300 53708 1352
rect 49148 1232 49200 1284
rect 51724 1232 51776 1284
rect 52368 1232 52420 1284
rect 50528 1164 50580 1216
rect 52920 1164 52972 1216
rect 54852 1300 54904 1352
rect 56324 1300 56376 1352
rect 54760 1232 54812 1284
rect 55680 1164 55732 1216
rect 59268 1343 59320 1352
rect 59268 1309 59277 1343
rect 59277 1309 59311 1343
rect 59311 1309 59320 1343
rect 59268 1300 59320 1309
rect 61200 1300 61252 1352
rect 62304 1300 62356 1352
rect 62580 1300 62632 1352
rect 63684 1343 63736 1352
rect 63684 1309 63693 1343
rect 63693 1309 63727 1343
rect 63727 1309 63736 1343
rect 63684 1300 63736 1309
rect 69940 1368 69992 1420
rect 66720 1300 66772 1352
rect 67640 1343 67692 1352
rect 67640 1309 67649 1343
rect 67649 1309 67683 1343
rect 67683 1309 67692 1343
rect 67640 1300 67692 1309
rect 68100 1300 68152 1352
rect 70584 1300 70636 1352
rect 70860 1300 70912 1352
rect 64604 1275 64656 1284
rect 64604 1241 64613 1275
rect 64613 1241 64647 1275
rect 64647 1241 64656 1275
rect 64604 1232 64656 1241
rect 65432 1232 65484 1284
rect 67548 1232 67600 1284
rect 72608 1232 72660 1284
rect 57336 1164 57388 1216
rect 65616 1164 65668 1216
rect 4210 1062 4262 1114
rect 4274 1062 4326 1114
rect 4338 1062 4390 1114
rect 4402 1062 4454 1114
rect 4466 1062 4518 1114
rect 14210 1062 14262 1114
rect 14274 1062 14326 1114
rect 14338 1062 14390 1114
rect 14402 1062 14454 1114
rect 14466 1062 14518 1114
rect 24210 1062 24262 1114
rect 24274 1062 24326 1114
rect 24338 1062 24390 1114
rect 24402 1062 24454 1114
rect 24466 1062 24518 1114
rect 34210 1062 34262 1114
rect 34274 1062 34326 1114
rect 34338 1062 34390 1114
rect 34402 1062 34454 1114
rect 34466 1062 34518 1114
rect 44210 1062 44262 1114
rect 44274 1062 44326 1114
rect 44338 1062 44390 1114
rect 44402 1062 44454 1114
rect 44466 1062 44518 1114
rect 54210 1062 54262 1114
rect 54274 1062 54326 1114
rect 54338 1062 54390 1114
rect 54402 1062 54454 1114
rect 54466 1062 54518 1114
rect 64210 1062 64262 1114
rect 64274 1062 64326 1114
rect 64338 1062 64390 1114
rect 64402 1062 64454 1114
rect 64466 1062 64518 1114
rect 74210 1062 74262 1114
rect 74274 1062 74326 1114
rect 74338 1062 74390 1114
rect 74402 1062 74454 1114
rect 74466 1062 74518 1114
rect 25688 960 25740 1012
rect 28264 960 28316 1012
rect 30840 960 30892 1012
rect 33324 960 33376 1012
rect 29828 892 29880 944
rect 34520 892 34572 944
rect 41420 960 41472 1012
rect 43904 960 43956 1012
rect 44088 960 44140 1012
rect 49148 960 49200 1012
rect 51724 960 51776 1012
rect 57336 960 57388 1012
rect 60280 960 60332 1012
rect 64604 960 64656 1012
rect 45192 892 45244 944
rect 48504 892 48556 944
rect 49608 892 49660 944
rect 27252 824 27304 876
rect 32588 824 32640 876
rect 33416 756 33468 808
rect 30932 688 30984 740
rect 47492 824 47544 876
rect 23112 76 23164 128
rect 65708 76 65760 128
<< metal2 >>
rect 71836 85434 72188 86000
rect 71836 85382 71858 85434
rect 71910 85382 71922 85434
rect 71974 85382 71986 85434
rect 72038 85382 72050 85434
rect 72102 85382 72114 85434
rect 72166 85382 72188 85434
rect 2112 84588 2216 84616
rect 2112 84532 2136 84588
rect 2192 84532 2216 84588
rect 2112 84508 2216 84532
rect 2112 84452 2136 84508
rect 2192 84452 2216 84508
rect 2112 84428 2216 84452
rect 2112 84372 2136 84428
rect 2192 84372 2216 84428
rect 2112 84348 2216 84372
rect 2112 84292 2136 84348
rect 2192 84292 2216 84348
rect 2112 84264 2216 84292
rect 5613 84588 5707 84616
rect 5613 84532 5632 84588
rect 5688 84532 5707 84588
rect 5613 84508 5707 84532
rect 5613 84452 5632 84508
rect 5688 84452 5707 84508
rect 5613 84428 5707 84452
rect 5613 84372 5632 84428
rect 5688 84372 5707 84428
rect 5613 84348 5707 84372
rect 5613 84292 5632 84348
rect 5688 84292 5707 84348
rect 5613 84264 5707 84292
rect 8503 84588 8597 84616
rect 8503 84532 8522 84588
rect 8578 84532 8597 84588
rect 8503 84508 8597 84532
rect 8503 84452 8522 84508
rect 8578 84452 8597 84508
rect 8503 84428 8597 84452
rect 8503 84372 8522 84428
rect 8578 84372 8597 84428
rect 8503 84348 8597 84372
rect 8503 84292 8522 84348
rect 8578 84292 8597 84348
rect 8503 84264 8597 84292
rect 11393 84588 11487 84616
rect 11393 84532 11412 84588
rect 11468 84532 11487 84588
rect 11393 84508 11487 84532
rect 11393 84452 11412 84508
rect 11468 84452 11487 84508
rect 11393 84428 11487 84452
rect 11393 84372 11412 84428
rect 11468 84372 11487 84428
rect 11393 84348 11487 84372
rect 11393 84292 11412 84348
rect 11468 84292 11487 84348
rect 11393 84264 11487 84292
rect 14283 84588 14377 84616
rect 14283 84532 14302 84588
rect 14358 84532 14377 84588
rect 14283 84508 14377 84532
rect 14283 84452 14302 84508
rect 14358 84452 14377 84508
rect 14283 84428 14377 84452
rect 14283 84372 14302 84428
rect 14358 84372 14377 84428
rect 14283 84348 14377 84372
rect 14283 84292 14302 84348
rect 14358 84292 14377 84348
rect 14283 84264 14377 84292
rect 17173 84588 17267 84616
rect 17173 84532 17192 84588
rect 17248 84532 17267 84588
rect 17173 84508 17267 84532
rect 17173 84452 17192 84508
rect 17248 84452 17267 84508
rect 17173 84428 17267 84452
rect 17173 84372 17192 84428
rect 17248 84372 17267 84428
rect 17173 84348 17267 84372
rect 17173 84292 17192 84348
rect 17248 84292 17267 84348
rect 17173 84264 17267 84292
rect 20063 84588 20157 84616
rect 20063 84532 20082 84588
rect 20138 84532 20157 84588
rect 20063 84508 20157 84532
rect 20063 84452 20082 84508
rect 20138 84452 20157 84508
rect 20063 84428 20157 84452
rect 20063 84372 20082 84428
rect 20138 84372 20157 84428
rect 20063 84348 20157 84372
rect 20063 84292 20082 84348
rect 20138 84292 20157 84348
rect 20063 84264 20157 84292
rect 22953 84588 23047 84616
rect 22953 84532 22972 84588
rect 23028 84532 23047 84588
rect 22953 84508 23047 84532
rect 22953 84452 22972 84508
rect 23028 84452 23047 84508
rect 22953 84428 23047 84452
rect 22953 84372 22972 84428
rect 23028 84372 23047 84428
rect 22953 84348 23047 84372
rect 22953 84292 22972 84348
rect 23028 84292 23047 84348
rect 22953 84264 23047 84292
rect 25843 84588 25937 84616
rect 25843 84532 25862 84588
rect 25918 84532 25937 84588
rect 25843 84508 25937 84532
rect 25843 84452 25862 84508
rect 25918 84452 25937 84508
rect 25843 84428 25937 84452
rect 25843 84372 25862 84428
rect 25918 84372 25937 84428
rect 25843 84348 25937 84372
rect 25843 84292 25862 84348
rect 25918 84292 25937 84348
rect 25843 84264 25937 84292
rect 28733 84588 28827 84616
rect 28733 84532 28752 84588
rect 28808 84532 28827 84588
rect 28733 84508 28827 84532
rect 28733 84452 28752 84508
rect 28808 84452 28827 84508
rect 28733 84428 28827 84452
rect 28733 84372 28752 84428
rect 28808 84372 28827 84428
rect 28733 84348 28827 84372
rect 28733 84292 28752 84348
rect 28808 84292 28827 84348
rect 28733 84264 28827 84292
rect 31623 84588 31717 84616
rect 31623 84532 31642 84588
rect 31698 84532 31717 84588
rect 31623 84508 31717 84532
rect 31623 84452 31642 84508
rect 31698 84452 31717 84508
rect 31623 84428 31717 84452
rect 31623 84372 31642 84428
rect 31698 84372 31717 84428
rect 31623 84348 31717 84372
rect 31623 84292 31642 84348
rect 31698 84292 31717 84348
rect 31623 84264 31717 84292
rect 34513 84588 34607 84616
rect 34513 84532 34532 84588
rect 34588 84532 34607 84588
rect 34513 84508 34607 84532
rect 34513 84452 34532 84508
rect 34588 84452 34607 84508
rect 34513 84428 34607 84452
rect 34513 84372 34532 84428
rect 34588 84372 34607 84428
rect 34513 84348 34607 84372
rect 34513 84292 34532 84348
rect 34588 84292 34607 84348
rect 34513 84264 34607 84292
rect 37403 84588 37497 84616
rect 37403 84532 37422 84588
rect 37478 84532 37497 84588
rect 37403 84508 37497 84532
rect 37403 84452 37422 84508
rect 37478 84452 37497 84508
rect 37403 84428 37497 84452
rect 37403 84372 37422 84428
rect 37478 84372 37497 84428
rect 37403 84348 37497 84372
rect 37403 84292 37422 84348
rect 37478 84292 37497 84348
rect 37403 84264 37497 84292
rect 40293 84588 40387 84616
rect 40293 84532 40312 84588
rect 40368 84532 40387 84588
rect 40293 84508 40387 84532
rect 40293 84452 40312 84508
rect 40368 84452 40387 84508
rect 40293 84428 40387 84452
rect 40293 84372 40312 84428
rect 40368 84372 40387 84428
rect 40293 84348 40387 84372
rect 40293 84292 40312 84348
rect 40368 84292 40387 84348
rect 40293 84264 40387 84292
rect 43183 84588 43277 84616
rect 43183 84532 43202 84588
rect 43258 84532 43277 84588
rect 43183 84508 43277 84532
rect 43183 84452 43202 84508
rect 43258 84452 43277 84508
rect 43183 84428 43277 84452
rect 43183 84372 43202 84428
rect 43258 84372 43277 84428
rect 43183 84348 43277 84372
rect 43183 84292 43202 84348
rect 43258 84292 43277 84348
rect 43183 84264 43277 84292
rect 46073 84588 46167 84616
rect 46073 84532 46092 84588
rect 46148 84532 46167 84588
rect 46073 84508 46167 84532
rect 46073 84452 46092 84508
rect 46148 84452 46167 84508
rect 46073 84428 46167 84452
rect 46073 84372 46092 84428
rect 46148 84372 46167 84428
rect 46073 84348 46167 84372
rect 46073 84292 46092 84348
rect 46148 84292 46167 84348
rect 46073 84264 46167 84292
rect 49081 84588 49175 84616
rect 49081 84532 49100 84588
rect 49156 84532 49175 84588
rect 49081 84508 49175 84532
rect 49081 84452 49100 84508
rect 49156 84452 49175 84508
rect 49081 84428 49175 84452
rect 49081 84372 49100 84428
rect 49156 84372 49175 84428
rect 49081 84348 49175 84372
rect 49081 84292 49100 84348
rect 49156 84292 49175 84348
rect 49081 84264 49175 84292
rect 52302 84588 52412 84616
rect 52302 84532 52329 84588
rect 52385 84532 52412 84588
rect 52302 84508 52412 84532
rect 52302 84452 52329 84508
rect 52385 84452 52412 84508
rect 52302 84428 52412 84452
rect 52302 84372 52329 84428
rect 52385 84372 52412 84428
rect 52302 84348 52412 84372
rect 52302 84292 52329 84348
rect 52385 84292 52412 84348
rect 52302 84264 52412 84292
rect 53694 84588 53822 84616
rect 53694 84532 53730 84588
rect 53786 84532 53822 84588
rect 53694 84508 53822 84532
rect 53694 84452 53730 84508
rect 53786 84452 53822 84508
rect 53694 84428 53822 84452
rect 53694 84372 53730 84428
rect 53786 84372 53822 84428
rect 53694 84348 53822 84372
rect 53694 84292 53730 84348
rect 53786 84292 53822 84348
rect 53694 84264 53822 84292
rect 53862 84588 53990 84616
rect 53862 84532 53898 84588
rect 53954 84532 53990 84588
rect 53862 84508 53990 84532
rect 53862 84452 53898 84508
rect 53954 84452 53990 84508
rect 53862 84428 53990 84452
rect 53862 84372 53898 84428
rect 53954 84372 53990 84428
rect 53862 84348 53990 84372
rect 53862 84292 53898 84348
rect 53954 84292 53990 84348
rect 53862 84264 53990 84292
rect 54606 84588 54734 84616
rect 54606 84532 54642 84588
rect 54698 84532 54734 84588
rect 54606 84508 54734 84532
rect 54606 84452 54642 84508
rect 54698 84452 54734 84508
rect 54606 84428 54734 84452
rect 54606 84372 54642 84428
rect 54698 84372 54734 84428
rect 54606 84348 54734 84372
rect 54606 84292 54642 84348
rect 54698 84292 54734 84348
rect 54606 84264 54734 84292
rect 55002 84588 55118 84616
rect 55002 84532 55032 84588
rect 55088 84532 55118 84588
rect 55002 84508 55118 84532
rect 55002 84452 55032 84508
rect 55088 84452 55118 84508
rect 55002 84428 55118 84452
rect 55002 84372 55032 84428
rect 55088 84372 55118 84428
rect 55002 84348 55118 84372
rect 55002 84292 55032 84348
rect 55088 84292 55118 84348
rect 55002 84264 55118 84292
rect 55712 84588 55840 84616
rect 55712 84532 55748 84588
rect 55804 84532 55840 84588
rect 55712 84508 55840 84532
rect 55712 84452 55748 84508
rect 55804 84452 55840 84508
rect 55712 84428 55840 84452
rect 55712 84372 55748 84428
rect 55804 84372 55840 84428
rect 55712 84348 55840 84372
rect 55712 84292 55748 84348
rect 55804 84292 55840 84348
rect 55712 84264 55840 84292
rect 56290 84588 56418 84616
rect 56290 84532 56326 84588
rect 56382 84532 56418 84588
rect 56290 84508 56418 84532
rect 56290 84452 56326 84508
rect 56382 84452 56418 84508
rect 56290 84428 56418 84452
rect 56290 84372 56326 84428
rect 56382 84372 56418 84428
rect 56290 84348 56418 84372
rect 56290 84292 56326 84348
rect 56382 84292 56418 84348
rect 56290 84264 56418 84292
rect 56741 84588 56857 84616
rect 56741 84532 56771 84588
rect 56827 84532 56857 84588
rect 56741 84508 56857 84532
rect 56741 84452 56771 84508
rect 56827 84452 56857 84508
rect 56741 84428 56857 84452
rect 56741 84372 56771 84428
rect 56827 84372 56857 84428
rect 56741 84348 56857 84372
rect 56741 84292 56771 84348
rect 56827 84292 56857 84348
rect 56741 84264 56857 84292
rect 57045 84588 57161 84616
rect 57045 84532 57075 84588
rect 57131 84532 57161 84588
rect 57045 84508 57161 84532
rect 57045 84452 57075 84508
rect 57131 84452 57161 84508
rect 57045 84428 57161 84452
rect 57045 84372 57075 84428
rect 57131 84372 57161 84428
rect 57045 84348 57161 84372
rect 57045 84292 57075 84348
rect 57131 84292 57161 84348
rect 57045 84264 57161 84292
rect 57887 84588 58003 84616
rect 57887 84532 57917 84588
rect 57973 84532 58003 84588
rect 57887 84508 58003 84532
rect 57887 84452 57917 84508
rect 57973 84452 58003 84508
rect 57887 84428 58003 84452
rect 57887 84372 57917 84428
rect 57973 84372 58003 84428
rect 57887 84348 58003 84372
rect 57887 84292 57917 84348
rect 57973 84292 58003 84348
rect 57887 84264 58003 84292
rect 58553 84588 58617 84616
rect 58553 84532 58557 84588
rect 58613 84532 58617 84588
rect 58553 84508 58617 84532
rect 58553 84452 58557 84508
rect 58613 84452 58617 84508
rect 58553 84428 58617 84452
rect 58553 84372 58557 84428
rect 58613 84372 58617 84428
rect 58553 84348 58617 84372
rect 58553 84292 58557 84348
rect 58613 84292 58617 84348
rect 58553 84264 58617 84292
rect 59110 84588 59226 84616
rect 59110 84532 59140 84588
rect 59196 84532 59226 84588
rect 59110 84508 59226 84532
rect 59110 84452 59140 84508
rect 59196 84452 59226 84508
rect 59110 84428 59226 84452
rect 59110 84372 59140 84428
rect 59196 84372 59226 84428
rect 59110 84348 59226 84372
rect 59110 84292 59140 84348
rect 59196 84292 59226 84348
rect 59110 84264 59226 84292
rect 60388 84588 60504 84616
rect 60388 84532 60418 84588
rect 60474 84532 60504 84588
rect 60388 84508 60504 84532
rect 60388 84452 60418 84508
rect 60474 84452 60504 84508
rect 60388 84428 60504 84452
rect 60388 84372 60418 84428
rect 60474 84372 60504 84428
rect 60388 84348 60504 84372
rect 60388 84292 60418 84348
rect 60474 84292 60504 84348
rect 60388 84264 60504 84292
rect 60546 84588 60662 84616
rect 60546 84532 60576 84588
rect 60632 84532 60662 84588
rect 60546 84508 60662 84532
rect 60546 84452 60576 84508
rect 60632 84452 60662 84508
rect 60546 84428 60662 84452
rect 60546 84372 60576 84428
rect 60632 84372 60662 84428
rect 60546 84348 60662 84372
rect 60546 84292 60576 84348
rect 60632 84292 60662 84348
rect 60546 84264 60662 84292
rect 62601 84588 62775 84616
rect 62601 84532 62620 84588
rect 62676 84532 62700 84588
rect 62756 84532 62775 84588
rect 62601 84508 62775 84532
rect 62601 84452 62620 84508
rect 62676 84452 62700 84508
rect 62756 84452 62775 84508
rect 62601 84428 62775 84452
rect 62601 84372 62620 84428
rect 62676 84372 62700 84428
rect 62756 84372 62775 84428
rect 62601 84348 62775 84372
rect 62601 84292 62620 84348
rect 62676 84292 62700 84348
rect 62756 84292 62775 84348
rect 62601 84264 62775 84292
rect 71836 84346 72188 85382
rect 71836 84294 71858 84346
rect 71910 84294 71922 84346
rect 71974 84294 71986 84346
rect 72038 84294 72050 84346
rect 72102 84294 72114 84346
rect 72166 84294 72188 84346
rect 63500 84244 63552 84250
rect 63500 84186 63552 84192
rect 63512 82414 63540 84186
rect 71836 83258 72188 84294
rect 71836 83206 71858 83258
rect 71910 83206 71922 83258
rect 71974 83206 71986 83258
rect 72038 83206 72050 83258
rect 72102 83206 72114 83258
rect 72166 83206 72188 83258
rect 66904 83156 66956 83162
rect 66904 83098 66956 83104
rect 63500 82408 63552 82414
rect 63500 82350 63552 82356
rect 2244 82236 2444 82264
rect 2244 82180 2276 82236
rect 2332 82180 2356 82236
rect 2412 82180 2444 82236
rect 2244 82156 2444 82180
rect 2244 82100 2276 82156
rect 2332 82100 2356 82156
rect 2412 82100 2444 82156
rect 2244 82076 2444 82100
rect 2244 82020 2276 82076
rect 2332 82020 2356 82076
rect 2412 82020 2444 82076
rect 2244 81996 2444 82020
rect 2244 81940 2276 81996
rect 2332 81940 2356 81996
rect 2412 81940 2444 81996
rect 2244 81912 2444 81940
rect 5466 82236 5560 82264
rect 5466 82180 5485 82236
rect 5541 82180 5560 82236
rect 5466 82156 5560 82180
rect 5466 82100 5485 82156
rect 5541 82100 5560 82156
rect 5466 82076 5560 82100
rect 5466 82020 5485 82076
rect 5541 82020 5560 82076
rect 5466 81996 5560 82020
rect 5466 81940 5485 81996
rect 5541 81940 5560 81996
rect 5466 81912 5560 81940
rect 8356 82236 8450 82264
rect 8356 82180 8375 82236
rect 8431 82180 8450 82236
rect 8356 82156 8450 82180
rect 8356 82100 8375 82156
rect 8431 82100 8450 82156
rect 8356 82076 8450 82100
rect 8356 82020 8375 82076
rect 8431 82020 8450 82076
rect 8356 81996 8450 82020
rect 8356 81940 8375 81996
rect 8431 81940 8450 81996
rect 8356 81912 8450 81940
rect 11246 82236 11340 82264
rect 11246 82180 11265 82236
rect 11321 82180 11340 82236
rect 11246 82156 11340 82180
rect 11246 82100 11265 82156
rect 11321 82100 11340 82156
rect 11246 82076 11340 82100
rect 11246 82020 11265 82076
rect 11321 82020 11340 82076
rect 11246 81996 11340 82020
rect 11246 81940 11265 81996
rect 11321 81940 11340 81996
rect 11246 81912 11340 81940
rect 14136 82236 14230 82264
rect 14136 82180 14155 82236
rect 14211 82180 14230 82236
rect 14136 82156 14230 82180
rect 14136 82100 14155 82156
rect 14211 82100 14230 82156
rect 14136 82076 14230 82100
rect 14136 82020 14155 82076
rect 14211 82020 14230 82076
rect 14136 81996 14230 82020
rect 14136 81940 14155 81996
rect 14211 81940 14230 81996
rect 14136 81912 14230 81940
rect 17026 82236 17120 82264
rect 17026 82180 17045 82236
rect 17101 82180 17120 82236
rect 17026 82156 17120 82180
rect 17026 82100 17045 82156
rect 17101 82100 17120 82156
rect 17026 82076 17120 82100
rect 17026 82020 17045 82076
rect 17101 82020 17120 82076
rect 17026 81996 17120 82020
rect 17026 81940 17045 81996
rect 17101 81940 17120 81996
rect 17026 81912 17120 81940
rect 19916 82236 20010 82264
rect 19916 82180 19935 82236
rect 19991 82180 20010 82236
rect 19916 82156 20010 82180
rect 19916 82100 19935 82156
rect 19991 82100 20010 82156
rect 19916 82076 20010 82100
rect 19916 82020 19935 82076
rect 19991 82020 20010 82076
rect 19916 81996 20010 82020
rect 19916 81940 19935 81996
rect 19991 81940 20010 81996
rect 19916 81912 20010 81940
rect 22806 82236 22900 82264
rect 22806 82180 22825 82236
rect 22881 82180 22900 82236
rect 22806 82156 22900 82180
rect 22806 82100 22825 82156
rect 22881 82100 22900 82156
rect 22806 82076 22900 82100
rect 22806 82020 22825 82076
rect 22881 82020 22900 82076
rect 22806 81996 22900 82020
rect 22806 81940 22825 81996
rect 22881 81940 22900 81996
rect 22806 81912 22900 81940
rect 25696 82236 25790 82264
rect 25696 82180 25715 82236
rect 25771 82180 25790 82236
rect 25696 82156 25790 82180
rect 25696 82100 25715 82156
rect 25771 82100 25790 82156
rect 25696 82076 25790 82100
rect 25696 82020 25715 82076
rect 25771 82020 25790 82076
rect 25696 81996 25790 82020
rect 25696 81940 25715 81996
rect 25771 81940 25790 81996
rect 25696 81912 25790 81940
rect 28586 82236 28680 82264
rect 28586 82180 28605 82236
rect 28661 82180 28680 82236
rect 28586 82156 28680 82180
rect 28586 82100 28605 82156
rect 28661 82100 28680 82156
rect 28586 82076 28680 82100
rect 28586 82020 28605 82076
rect 28661 82020 28680 82076
rect 28586 81996 28680 82020
rect 28586 81940 28605 81996
rect 28661 81940 28680 81996
rect 28586 81912 28680 81940
rect 31476 82236 31570 82264
rect 31476 82180 31495 82236
rect 31551 82180 31570 82236
rect 31476 82156 31570 82180
rect 31476 82100 31495 82156
rect 31551 82100 31570 82156
rect 31476 82076 31570 82100
rect 31476 82020 31495 82076
rect 31551 82020 31570 82076
rect 31476 81996 31570 82020
rect 31476 81940 31495 81996
rect 31551 81940 31570 81996
rect 31476 81912 31570 81940
rect 34366 82236 34460 82264
rect 34366 82180 34385 82236
rect 34441 82180 34460 82236
rect 34366 82156 34460 82180
rect 34366 82100 34385 82156
rect 34441 82100 34460 82156
rect 34366 82076 34460 82100
rect 34366 82020 34385 82076
rect 34441 82020 34460 82076
rect 34366 81996 34460 82020
rect 34366 81940 34385 81996
rect 34441 81940 34460 81996
rect 34366 81912 34460 81940
rect 37256 82236 37350 82264
rect 37256 82180 37275 82236
rect 37331 82180 37350 82236
rect 37256 82156 37350 82180
rect 37256 82100 37275 82156
rect 37331 82100 37350 82156
rect 37256 82076 37350 82100
rect 37256 82020 37275 82076
rect 37331 82020 37350 82076
rect 37256 81996 37350 82020
rect 37256 81940 37275 81996
rect 37331 81940 37350 81996
rect 37256 81912 37350 81940
rect 40146 82236 40240 82264
rect 40146 82180 40165 82236
rect 40221 82180 40240 82236
rect 40146 82156 40240 82180
rect 40146 82100 40165 82156
rect 40221 82100 40240 82156
rect 40146 82076 40240 82100
rect 40146 82020 40165 82076
rect 40221 82020 40240 82076
rect 40146 81996 40240 82020
rect 40146 81940 40165 81996
rect 40221 81940 40240 81996
rect 40146 81912 40240 81940
rect 43036 82236 43130 82264
rect 43036 82180 43055 82236
rect 43111 82180 43130 82236
rect 43036 82156 43130 82180
rect 43036 82100 43055 82156
rect 43111 82100 43130 82156
rect 43036 82076 43130 82100
rect 43036 82020 43055 82076
rect 43111 82020 43130 82076
rect 43036 81996 43130 82020
rect 43036 81940 43055 81996
rect 43111 81940 43130 81996
rect 43036 81912 43130 81940
rect 45926 82236 46020 82264
rect 45926 82180 45945 82236
rect 46001 82180 46020 82236
rect 45926 82156 46020 82180
rect 45926 82100 45945 82156
rect 46001 82100 46020 82156
rect 45926 82076 46020 82100
rect 45926 82020 45945 82076
rect 46001 82020 46020 82076
rect 45926 81996 46020 82020
rect 45926 81940 45945 81996
rect 46001 81940 46020 81996
rect 45926 81912 46020 81940
rect 48873 82236 48967 82264
rect 48873 82180 48892 82236
rect 48948 82180 48967 82236
rect 48873 82156 48967 82180
rect 48873 82100 48892 82156
rect 48948 82100 48967 82156
rect 48873 82076 48967 82100
rect 48873 82020 48892 82076
rect 48948 82020 48967 82076
rect 48873 81996 48967 82020
rect 48873 81940 48892 81996
rect 48948 81940 48967 81996
rect 48873 81912 48967 81940
rect 49722 82236 49922 82264
rect 49722 82180 49754 82236
rect 49810 82180 49834 82236
rect 49890 82180 49922 82236
rect 49722 82156 49922 82180
rect 49722 82100 49754 82156
rect 49810 82100 49834 82156
rect 49890 82100 49922 82156
rect 49722 82076 49922 82100
rect 49722 82020 49754 82076
rect 49810 82020 49834 82076
rect 49890 82020 49922 82076
rect 49722 81996 49922 82020
rect 49722 81940 49754 81996
rect 49810 81940 49834 81996
rect 49890 81940 49922 81996
rect 49722 81912 49922 81940
rect 53012 82236 53140 82264
rect 53012 82180 53048 82236
rect 53104 82180 53140 82236
rect 53012 82156 53140 82180
rect 53012 82100 53048 82156
rect 53104 82100 53140 82156
rect 53012 82076 53140 82100
rect 53012 82020 53048 82076
rect 53104 82020 53140 82076
rect 53012 81996 53140 82020
rect 53012 81940 53048 81996
rect 53104 81940 53140 81996
rect 53012 81912 53140 81940
rect 53170 82236 53298 82264
rect 53170 82180 53206 82236
rect 53262 82180 53298 82236
rect 53170 82156 53298 82180
rect 53170 82100 53206 82156
rect 53262 82100 53298 82156
rect 53170 82076 53298 82100
rect 53170 82020 53206 82076
rect 53262 82020 53298 82076
rect 53170 81996 53298 82020
rect 53170 81940 53206 81996
rect 53262 81940 53298 81996
rect 53170 81912 53298 81940
rect 53526 82236 53654 82264
rect 53526 82180 53562 82236
rect 53618 82180 53654 82236
rect 53526 82156 53654 82180
rect 53526 82100 53562 82156
rect 53618 82100 53654 82156
rect 53526 82076 53654 82100
rect 53526 82020 53562 82076
rect 53618 82020 53654 82076
rect 53526 81996 53654 82020
rect 53526 81940 53562 81996
rect 53618 81940 53654 81996
rect 53526 81912 53654 81940
rect 54844 82236 54972 82264
rect 54844 82180 54880 82236
rect 54936 82180 54972 82236
rect 54844 82156 54972 82180
rect 54844 82100 54880 82156
rect 54936 82100 54972 82156
rect 54844 82076 54972 82100
rect 54844 82020 54880 82076
rect 54936 82020 54972 82076
rect 54844 81996 54972 82020
rect 54844 81940 54880 81996
rect 54936 81940 54972 81996
rect 54844 81912 54972 81940
rect 55437 82236 55565 82264
rect 55437 82180 55473 82236
rect 55529 82180 55565 82236
rect 55437 82156 55565 82180
rect 55437 82100 55473 82156
rect 55529 82100 55565 82156
rect 55437 82076 55565 82100
rect 55437 82020 55473 82076
rect 55529 82020 55565 82076
rect 55437 81996 55565 82020
rect 55437 81940 55473 81996
rect 55529 81940 55565 81996
rect 55437 81912 55565 81940
rect 56583 82236 56711 82264
rect 56583 82180 56619 82236
rect 56675 82180 56711 82236
rect 56583 82156 56711 82180
rect 56583 82100 56619 82156
rect 56675 82100 56711 82156
rect 56583 82076 56711 82100
rect 56583 82020 56619 82076
rect 56675 82020 56711 82076
rect 56583 81996 56711 82020
rect 56583 81940 56619 81996
rect 56675 81940 56711 81996
rect 56583 81912 56711 81940
rect 58033 82236 58213 82264
rect 58033 82180 58055 82236
rect 58111 82180 58135 82236
rect 58191 82180 58213 82236
rect 58033 82156 58213 82180
rect 58033 82100 58055 82156
rect 58111 82100 58135 82156
rect 58191 82100 58213 82156
rect 58033 82076 58213 82100
rect 58033 82020 58055 82076
rect 58111 82020 58135 82076
rect 58191 82020 58213 82076
rect 58033 81996 58213 82020
rect 58033 81940 58055 81996
rect 58111 81940 58135 81996
rect 58191 81940 58213 81996
rect 58033 81912 58213 81940
rect 59256 82236 59396 82264
rect 59256 82180 59298 82236
rect 59354 82180 59396 82236
rect 59256 82156 59396 82180
rect 59256 82100 59298 82156
rect 59354 82100 59396 82156
rect 59256 82076 59396 82100
rect 59256 82020 59298 82076
rect 59354 82020 59396 82076
rect 59256 81996 59396 82020
rect 59256 81940 59298 81996
rect 59354 81940 59396 81996
rect 59256 81912 59396 81940
rect 59426 82236 59542 82264
rect 59426 82180 59456 82236
rect 59512 82180 59542 82236
rect 59426 82156 59542 82180
rect 59426 82100 59456 82156
rect 59512 82100 59542 82156
rect 59426 82076 59542 82100
rect 59426 82020 59456 82076
rect 59512 82020 59542 82076
rect 59426 81996 59542 82020
rect 59426 81940 59456 81996
rect 59512 81940 59542 81996
rect 59426 81912 59542 81940
rect 59734 82236 59850 82264
rect 59734 82180 59764 82236
rect 59820 82180 59850 82236
rect 59734 82156 59850 82180
rect 59734 82100 59764 82156
rect 59820 82100 59850 82156
rect 59734 82076 59850 82100
rect 59734 82020 59764 82076
rect 59820 82020 59850 82076
rect 59734 81996 59850 82020
rect 59734 81940 59764 81996
rect 59820 81940 59850 81996
rect 59734 81912 59850 81940
rect 59880 82236 59996 82264
rect 59880 82180 59910 82236
rect 59966 82180 59996 82236
rect 59880 82156 59996 82180
rect 59880 82100 59910 82156
rect 59966 82100 59996 82156
rect 59880 82076 59996 82100
rect 59880 82020 59910 82076
rect 59966 82020 59996 82076
rect 59880 81996 59996 82020
rect 59880 81940 59910 81996
rect 59966 81940 59996 81996
rect 59880 81912 59996 81940
rect 60026 82236 60202 82264
rect 60026 82180 60046 82236
rect 60102 82180 60126 82236
rect 60182 82180 60202 82236
rect 60026 82156 60202 82180
rect 60026 82100 60046 82156
rect 60102 82100 60126 82156
rect 60182 82100 60202 82156
rect 60026 82076 60202 82100
rect 60026 82020 60046 82076
rect 60102 82020 60126 82076
rect 60182 82020 60202 82076
rect 60026 81996 60202 82020
rect 60026 81940 60046 81996
rect 60102 81940 60126 81996
rect 60182 81940 60202 81996
rect 60026 81912 60202 81940
rect 62399 82236 62573 82264
rect 62399 82180 62418 82236
rect 62474 82180 62498 82236
rect 62554 82180 62573 82236
rect 62399 82156 62573 82180
rect 62399 82100 62418 82156
rect 62474 82100 62498 82156
rect 62554 82100 62573 82156
rect 62399 82076 62573 82100
rect 62399 82020 62418 82076
rect 62474 82020 62498 82076
rect 62554 82020 62573 82076
rect 62399 81996 62573 82020
rect 62399 81940 62418 81996
rect 62474 81940 62498 81996
rect 62554 81940 62573 81996
rect 62399 81912 62573 81940
rect 63512 80034 63540 82350
rect 66720 80980 66772 80986
rect 66720 80922 66772 80928
rect 63500 80028 63552 80034
rect 63500 79970 63552 79976
rect 63512 78062 63540 79970
rect 65616 78736 65668 78742
rect 65616 78678 65668 78684
rect 63500 78056 63552 78062
rect 63500 77998 63552 78004
rect 63592 77444 63644 77450
rect 63592 77386 63644 77392
rect 63500 76742 63552 76748
rect 63500 76684 63552 76690
rect 2112 74588 2216 74616
rect 2112 74532 2136 74588
rect 2192 74532 2216 74588
rect 2112 74508 2216 74532
rect 2112 74452 2136 74508
rect 2192 74452 2216 74508
rect 2112 74428 2216 74452
rect 2112 74372 2136 74428
rect 2192 74372 2216 74428
rect 2112 74348 2216 74372
rect 2112 74292 2136 74348
rect 2192 74292 2216 74348
rect 2112 74264 2216 74292
rect 5613 74588 5707 74616
rect 5613 74532 5632 74588
rect 5688 74532 5707 74588
rect 5613 74508 5707 74532
rect 5613 74452 5632 74508
rect 5688 74452 5707 74508
rect 5613 74428 5707 74452
rect 5613 74372 5632 74428
rect 5688 74372 5707 74428
rect 5613 74348 5707 74372
rect 5613 74292 5632 74348
rect 5688 74292 5707 74348
rect 5613 74264 5707 74292
rect 8503 74588 8597 74616
rect 8503 74532 8522 74588
rect 8578 74532 8597 74588
rect 8503 74508 8597 74532
rect 8503 74452 8522 74508
rect 8578 74452 8597 74508
rect 8503 74428 8597 74452
rect 8503 74372 8522 74428
rect 8578 74372 8597 74428
rect 8503 74348 8597 74372
rect 8503 74292 8522 74348
rect 8578 74292 8597 74348
rect 8503 74264 8597 74292
rect 11393 74588 11487 74616
rect 11393 74532 11412 74588
rect 11468 74532 11487 74588
rect 11393 74508 11487 74532
rect 11393 74452 11412 74508
rect 11468 74452 11487 74508
rect 11393 74428 11487 74452
rect 11393 74372 11412 74428
rect 11468 74372 11487 74428
rect 11393 74348 11487 74372
rect 11393 74292 11412 74348
rect 11468 74292 11487 74348
rect 11393 74264 11487 74292
rect 14283 74588 14377 74616
rect 14283 74532 14302 74588
rect 14358 74532 14377 74588
rect 14283 74508 14377 74532
rect 14283 74452 14302 74508
rect 14358 74452 14377 74508
rect 14283 74428 14377 74452
rect 14283 74372 14302 74428
rect 14358 74372 14377 74428
rect 14283 74348 14377 74372
rect 14283 74292 14302 74348
rect 14358 74292 14377 74348
rect 14283 74264 14377 74292
rect 17173 74588 17267 74616
rect 17173 74532 17192 74588
rect 17248 74532 17267 74588
rect 17173 74508 17267 74532
rect 17173 74452 17192 74508
rect 17248 74452 17267 74508
rect 17173 74428 17267 74452
rect 17173 74372 17192 74428
rect 17248 74372 17267 74428
rect 17173 74348 17267 74372
rect 17173 74292 17192 74348
rect 17248 74292 17267 74348
rect 17173 74264 17267 74292
rect 20063 74588 20157 74616
rect 20063 74532 20082 74588
rect 20138 74532 20157 74588
rect 20063 74508 20157 74532
rect 20063 74452 20082 74508
rect 20138 74452 20157 74508
rect 20063 74428 20157 74452
rect 20063 74372 20082 74428
rect 20138 74372 20157 74428
rect 20063 74348 20157 74372
rect 20063 74292 20082 74348
rect 20138 74292 20157 74348
rect 20063 74264 20157 74292
rect 22953 74588 23047 74616
rect 22953 74532 22972 74588
rect 23028 74532 23047 74588
rect 22953 74508 23047 74532
rect 22953 74452 22972 74508
rect 23028 74452 23047 74508
rect 22953 74428 23047 74452
rect 22953 74372 22972 74428
rect 23028 74372 23047 74428
rect 22953 74348 23047 74372
rect 22953 74292 22972 74348
rect 23028 74292 23047 74348
rect 22953 74264 23047 74292
rect 25843 74588 25937 74616
rect 25843 74532 25862 74588
rect 25918 74532 25937 74588
rect 25843 74508 25937 74532
rect 25843 74452 25862 74508
rect 25918 74452 25937 74508
rect 25843 74428 25937 74452
rect 25843 74372 25862 74428
rect 25918 74372 25937 74428
rect 25843 74348 25937 74372
rect 25843 74292 25862 74348
rect 25918 74292 25937 74348
rect 25843 74264 25937 74292
rect 28733 74588 28827 74616
rect 28733 74532 28752 74588
rect 28808 74532 28827 74588
rect 28733 74508 28827 74532
rect 28733 74452 28752 74508
rect 28808 74452 28827 74508
rect 28733 74428 28827 74452
rect 28733 74372 28752 74428
rect 28808 74372 28827 74428
rect 28733 74348 28827 74372
rect 28733 74292 28752 74348
rect 28808 74292 28827 74348
rect 28733 74264 28827 74292
rect 31623 74588 31717 74616
rect 31623 74532 31642 74588
rect 31698 74532 31717 74588
rect 31623 74508 31717 74532
rect 31623 74452 31642 74508
rect 31698 74452 31717 74508
rect 31623 74428 31717 74452
rect 31623 74372 31642 74428
rect 31698 74372 31717 74428
rect 31623 74348 31717 74372
rect 31623 74292 31642 74348
rect 31698 74292 31717 74348
rect 31623 74264 31717 74292
rect 34513 74588 34607 74616
rect 34513 74532 34532 74588
rect 34588 74532 34607 74588
rect 34513 74508 34607 74532
rect 34513 74452 34532 74508
rect 34588 74452 34607 74508
rect 34513 74428 34607 74452
rect 34513 74372 34532 74428
rect 34588 74372 34607 74428
rect 34513 74348 34607 74372
rect 34513 74292 34532 74348
rect 34588 74292 34607 74348
rect 34513 74264 34607 74292
rect 37403 74588 37497 74616
rect 37403 74532 37422 74588
rect 37478 74532 37497 74588
rect 37403 74508 37497 74532
rect 37403 74452 37422 74508
rect 37478 74452 37497 74508
rect 37403 74428 37497 74452
rect 37403 74372 37422 74428
rect 37478 74372 37497 74428
rect 37403 74348 37497 74372
rect 37403 74292 37422 74348
rect 37478 74292 37497 74348
rect 37403 74264 37497 74292
rect 40293 74588 40387 74616
rect 40293 74532 40312 74588
rect 40368 74532 40387 74588
rect 40293 74508 40387 74532
rect 40293 74452 40312 74508
rect 40368 74452 40387 74508
rect 40293 74428 40387 74452
rect 40293 74372 40312 74428
rect 40368 74372 40387 74428
rect 40293 74348 40387 74372
rect 40293 74292 40312 74348
rect 40368 74292 40387 74348
rect 40293 74264 40387 74292
rect 43183 74588 43277 74616
rect 43183 74532 43202 74588
rect 43258 74532 43277 74588
rect 43183 74508 43277 74532
rect 43183 74452 43202 74508
rect 43258 74452 43277 74508
rect 43183 74428 43277 74452
rect 43183 74372 43202 74428
rect 43258 74372 43277 74428
rect 43183 74348 43277 74372
rect 43183 74292 43202 74348
rect 43258 74292 43277 74348
rect 43183 74264 43277 74292
rect 46073 74588 46167 74616
rect 46073 74532 46092 74588
rect 46148 74532 46167 74588
rect 46073 74508 46167 74532
rect 46073 74452 46092 74508
rect 46148 74452 46167 74508
rect 46073 74428 46167 74452
rect 46073 74372 46092 74428
rect 46148 74372 46167 74428
rect 46073 74348 46167 74372
rect 46073 74292 46092 74348
rect 46148 74292 46167 74348
rect 46073 74264 46167 74292
rect 49081 74588 49175 74616
rect 49081 74532 49100 74588
rect 49156 74532 49175 74588
rect 49081 74508 49175 74532
rect 49081 74452 49100 74508
rect 49156 74452 49175 74508
rect 49081 74428 49175 74452
rect 49081 74372 49100 74428
rect 49156 74372 49175 74428
rect 49081 74348 49175 74372
rect 49081 74292 49100 74348
rect 49156 74292 49175 74348
rect 49081 74264 49175 74292
rect 52302 74588 52412 74616
rect 52302 74532 52329 74588
rect 52385 74532 52412 74588
rect 52302 74508 52412 74532
rect 52302 74452 52329 74508
rect 52385 74452 52412 74508
rect 52302 74428 52412 74452
rect 52302 74372 52329 74428
rect 52385 74372 52412 74428
rect 52302 74348 52412 74372
rect 52302 74292 52329 74348
rect 52385 74292 52412 74348
rect 52302 74264 52412 74292
rect 53694 74588 53822 74616
rect 53694 74532 53730 74588
rect 53786 74532 53822 74588
rect 53694 74508 53822 74532
rect 53694 74452 53730 74508
rect 53786 74452 53822 74508
rect 53694 74428 53822 74452
rect 53694 74372 53730 74428
rect 53786 74372 53822 74428
rect 53694 74348 53822 74372
rect 53694 74292 53730 74348
rect 53786 74292 53822 74348
rect 53694 74264 53822 74292
rect 53862 74588 53990 74616
rect 53862 74532 53898 74588
rect 53954 74532 53990 74588
rect 53862 74508 53990 74532
rect 53862 74452 53898 74508
rect 53954 74452 53990 74508
rect 53862 74428 53990 74452
rect 53862 74372 53898 74428
rect 53954 74372 53990 74428
rect 53862 74348 53990 74372
rect 53862 74292 53898 74348
rect 53954 74292 53990 74348
rect 53862 74264 53990 74292
rect 54606 74588 54734 74616
rect 54606 74532 54642 74588
rect 54698 74532 54734 74588
rect 54606 74508 54734 74532
rect 54606 74452 54642 74508
rect 54698 74452 54734 74508
rect 54606 74428 54734 74452
rect 54606 74372 54642 74428
rect 54698 74372 54734 74428
rect 54606 74348 54734 74372
rect 54606 74292 54642 74348
rect 54698 74292 54734 74348
rect 54606 74264 54734 74292
rect 55002 74588 55118 74616
rect 55002 74532 55032 74588
rect 55088 74532 55118 74588
rect 55002 74508 55118 74532
rect 55002 74452 55032 74508
rect 55088 74452 55118 74508
rect 55002 74428 55118 74452
rect 55002 74372 55032 74428
rect 55088 74372 55118 74428
rect 55002 74348 55118 74372
rect 55002 74292 55032 74348
rect 55088 74292 55118 74348
rect 55002 74264 55118 74292
rect 55712 74588 55840 74616
rect 55712 74532 55748 74588
rect 55804 74532 55840 74588
rect 55712 74508 55840 74532
rect 55712 74452 55748 74508
rect 55804 74452 55840 74508
rect 55712 74428 55840 74452
rect 55712 74372 55748 74428
rect 55804 74372 55840 74428
rect 55712 74348 55840 74372
rect 55712 74292 55748 74348
rect 55804 74292 55840 74348
rect 55712 74264 55840 74292
rect 56290 74588 56418 74616
rect 56290 74532 56326 74588
rect 56382 74532 56418 74588
rect 56290 74508 56418 74532
rect 56290 74452 56326 74508
rect 56382 74452 56418 74508
rect 56290 74428 56418 74452
rect 56290 74372 56326 74428
rect 56382 74372 56418 74428
rect 56290 74348 56418 74372
rect 56290 74292 56326 74348
rect 56382 74292 56418 74348
rect 56290 74264 56418 74292
rect 56741 74588 56857 74616
rect 56741 74532 56771 74588
rect 56827 74532 56857 74588
rect 56741 74508 56857 74532
rect 56741 74452 56771 74508
rect 56827 74452 56857 74508
rect 56741 74428 56857 74452
rect 56741 74372 56771 74428
rect 56827 74372 56857 74428
rect 56741 74348 56857 74372
rect 56741 74292 56771 74348
rect 56827 74292 56857 74348
rect 56741 74264 56857 74292
rect 57045 74588 57161 74616
rect 57045 74532 57075 74588
rect 57131 74532 57161 74588
rect 57045 74508 57161 74532
rect 57045 74452 57075 74508
rect 57131 74452 57161 74508
rect 57045 74428 57161 74452
rect 57045 74372 57075 74428
rect 57131 74372 57161 74428
rect 57045 74348 57161 74372
rect 57045 74292 57075 74348
rect 57131 74292 57161 74348
rect 57045 74264 57161 74292
rect 57887 74588 58003 74616
rect 57887 74532 57917 74588
rect 57973 74532 58003 74588
rect 57887 74508 58003 74532
rect 57887 74452 57917 74508
rect 57973 74452 58003 74508
rect 57887 74428 58003 74452
rect 57887 74372 57917 74428
rect 57973 74372 58003 74428
rect 57887 74348 58003 74372
rect 57887 74292 57917 74348
rect 57973 74292 58003 74348
rect 57887 74264 58003 74292
rect 58553 74588 58617 74616
rect 58553 74532 58557 74588
rect 58613 74532 58617 74588
rect 58553 74508 58617 74532
rect 58553 74452 58557 74508
rect 58613 74452 58617 74508
rect 58553 74428 58617 74452
rect 58553 74372 58557 74428
rect 58613 74372 58617 74428
rect 58553 74348 58617 74372
rect 58553 74292 58557 74348
rect 58613 74292 58617 74348
rect 58553 74264 58617 74292
rect 59110 74588 59226 74616
rect 59110 74532 59140 74588
rect 59196 74532 59226 74588
rect 59110 74508 59226 74532
rect 59110 74452 59140 74508
rect 59196 74452 59226 74508
rect 59110 74428 59226 74452
rect 59110 74372 59140 74428
rect 59196 74372 59226 74428
rect 59110 74348 59226 74372
rect 59110 74292 59140 74348
rect 59196 74292 59226 74348
rect 59110 74264 59226 74292
rect 60388 74588 60504 74616
rect 60388 74532 60418 74588
rect 60474 74532 60504 74588
rect 60388 74508 60504 74532
rect 60388 74452 60418 74508
rect 60474 74452 60504 74508
rect 60388 74428 60504 74452
rect 60388 74372 60418 74428
rect 60474 74372 60504 74428
rect 60388 74348 60504 74372
rect 60388 74292 60418 74348
rect 60474 74292 60504 74348
rect 60388 74264 60504 74292
rect 60546 74588 60662 74616
rect 60546 74532 60576 74588
rect 60632 74532 60662 74588
rect 60546 74508 60662 74532
rect 60546 74452 60576 74508
rect 60632 74452 60662 74508
rect 60546 74428 60662 74452
rect 60546 74372 60576 74428
rect 60632 74372 60662 74428
rect 60546 74348 60662 74372
rect 60546 74292 60576 74348
rect 60632 74292 60662 74348
rect 60546 74264 60662 74292
rect 62601 74588 62775 74616
rect 62601 74532 62620 74588
rect 62676 74532 62700 74588
rect 62756 74532 62775 74588
rect 62601 74508 62775 74532
rect 62601 74452 62620 74508
rect 62676 74452 62700 74508
rect 62756 74452 62775 74508
rect 62601 74428 62775 74452
rect 62601 74372 62620 74428
rect 62676 74372 62700 74428
rect 62756 74372 62775 74428
rect 62601 74348 62775 74372
rect 62601 74292 62620 74348
rect 62676 74292 62700 74348
rect 62756 74292 62775 74348
rect 62601 74264 62775 74292
rect 2244 72236 2444 72264
rect 2244 72180 2276 72236
rect 2332 72180 2356 72236
rect 2412 72180 2444 72236
rect 2244 72156 2444 72180
rect 2244 72100 2276 72156
rect 2332 72100 2356 72156
rect 2412 72100 2444 72156
rect 2244 72076 2444 72100
rect 2244 72020 2276 72076
rect 2332 72020 2356 72076
rect 2412 72020 2444 72076
rect 2244 71996 2444 72020
rect 2244 71940 2276 71996
rect 2332 71940 2356 71996
rect 2412 71940 2444 71996
rect 2244 71912 2444 71940
rect 5466 72236 5560 72264
rect 5466 72180 5485 72236
rect 5541 72180 5560 72236
rect 5466 72156 5560 72180
rect 5466 72100 5485 72156
rect 5541 72100 5560 72156
rect 5466 72076 5560 72100
rect 5466 72020 5485 72076
rect 5541 72020 5560 72076
rect 5466 71996 5560 72020
rect 5466 71940 5485 71996
rect 5541 71940 5560 71996
rect 5466 71912 5560 71940
rect 8356 72236 8450 72264
rect 8356 72180 8375 72236
rect 8431 72180 8450 72236
rect 8356 72156 8450 72180
rect 8356 72100 8375 72156
rect 8431 72100 8450 72156
rect 8356 72076 8450 72100
rect 8356 72020 8375 72076
rect 8431 72020 8450 72076
rect 8356 71996 8450 72020
rect 8356 71940 8375 71996
rect 8431 71940 8450 71996
rect 8356 71912 8450 71940
rect 11246 72236 11340 72264
rect 11246 72180 11265 72236
rect 11321 72180 11340 72236
rect 11246 72156 11340 72180
rect 11246 72100 11265 72156
rect 11321 72100 11340 72156
rect 11246 72076 11340 72100
rect 11246 72020 11265 72076
rect 11321 72020 11340 72076
rect 11246 71996 11340 72020
rect 11246 71940 11265 71996
rect 11321 71940 11340 71996
rect 11246 71912 11340 71940
rect 14136 72236 14230 72264
rect 14136 72180 14155 72236
rect 14211 72180 14230 72236
rect 14136 72156 14230 72180
rect 14136 72100 14155 72156
rect 14211 72100 14230 72156
rect 14136 72076 14230 72100
rect 14136 72020 14155 72076
rect 14211 72020 14230 72076
rect 14136 71996 14230 72020
rect 14136 71940 14155 71996
rect 14211 71940 14230 71996
rect 14136 71912 14230 71940
rect 17026 72236 17120 72264
rect 17026 72180 17045 72236
rect 17101 72180 17120 72236
rect 17026 72156 17120 72180
rect 17026 72100 17045 72156
rect 17101 72100 17120 72156
rect 17026 72076 17120 72100
rect 17026 72020 17045 72076
rect 17101 72020 17120 72076
rect 17026 71996 17120 72020
rect 17026 71940 17045 71996
rect 17101 71940 17120 71996
rect 17026 71912 17120 71940
rect 19916 72236 20010 72264
rect 19916 72180 19935 72236
rect 19991 72180 20010 72236
rect 19916 72156 20010 72180
rect 19916 72100 19935 72156
rect 19991 72100 20010 72156
rect 19916 72076 20010 72100
rect 19916 72020 19935 72076
rect 19991 72020 20010 72076
rect 19916 71996 20010 72020
rect 19916 71940 19935 71996
rect 19991 71940 20010 71996
rect 19916 71912 20010 71940
rect 22806 72236 22900 72264
rect 22806 72180 22825 72236
rect 22881 72180 22900 72236
rect 22806 72156 22900 72180
rect 22806 72100 22825 72156
rect 22881 72100 22900 72156
rect 22806 72076 22900 72100
rect 22806 72020 22825 72076
rect 22881 72020 22900 72076
rect 22806 71996 22900 72020
rect 22806 71940 22825 71996
rect 22881 71940 22900 71996
rect 22806 71912 22900 71940
rect 25696 72236 25790 72264
rect 25696 72180 25715 72236
rect 25771 72180 25790 72236
rect 25696 72156 25790 72180
rect 25696 72100 25715 72156
rect 25771 72100 25790 72156
rect 25696 72076 25790 72100
rect 25696 72020 25715 72076
rect 25771 72020 25790 72076
rect 25696 71996 25790 72020
rect 25696 71940 25715 71996
rect 25771 71940 25790 71996
rect 25696 71912 25790 71940
rect 28586 72236 28680 72264
rect 28586 72180 28605 72236
rect 28661 72180 28680 72236
rect 28586 72156 28680 72180
rect 28586 72100 28605 72156
rect 28661 72100 28680 72156
rect 28586 72076 28680 72100
rect 28586 72020 28605 72076
rect 28661 72020 28680 72076
rect 28586 71996 28680 72020
rect 28586 71940 28605 71996
rect 28661 71940 28680 71996
rect 28586 71912 28680 71940
rect 31476 72236 31570 72264
rect 31476 72180 31495 72236
rect 31551 72180 31570 72236
rect 31476 72156 31570 72180
rect 31476 72100 31495 72156
rect 31551 72100 31570 72156
rect 31476 72076 31570 72100
rect 31476 72020 31495 72076
rect 31551 72020 31570 72076
rect 31476 71996 31570 72020
rect 31476 71940 31495 71996
rect 31551 71940 31570 71996
rect 31476 71912 31570 71940
rect 34366 72236 34460 72264
rect 34366 72180 34385 72236
rect 34441 72180 34460 72236
rect 34366 72156 34460 72180
rect 34366 72100 34385 72156
rect 34441 72100 34460 72156
rect 34366 72076 34460 72100
rect 34366 72020 34385 72076
rect 34441 72020 34460 72076
rect 34366 71996 34460 72020
rect 34366 71940 34385 71996
rect 34441 71940 34460 71996
rect 34366 71912 34460 71940
rect 37256 72236 37350 72264
rect 37256 72180 37275 72236
rect 37331 72180 37350 72236
rect 37256 72156 37350 72180
rect 37256 72100 37275 72156
rect 37331 72100 37350 72156
rect 37256 72076 37350 72100
rect 37256 72020 37275 72076
rect 37331 72020 37350 72076
rect 37256 71996 37350 72020
rect 37256 71940 37275 71996
rect 37331 71940 37350 71996
rect 37256 71912 37350 71940
rect 40146 72236 40240 72264
rect 40146 72180 40165 72236
rect 40221 72180 40240 72236
rect 40146 72156 40240 72180
rect 40146 72100 40165 72156
rect 40221 72100 40240 72156
rect 40146 72076 40240 72100
rect 40146 72020 40165 72076
rect 40221 72020 40240 72076
rect 40146 71996 40240 72020
rect 40146 71940 40165 71996
rect 40221 71940 40240 71996
rect 40146 71912 40240 71940
rect 43036 72236 43130 72264
rect 43036 72180 43055 72236
rect 43111 72180 43130 72236
rect 43036 72156 43130 72180
rect 43036 72100 43055 72156
rect 43111 72100 43130 72156
rect 43036 72076 43130 72100
rect 43036 72020 43055 72076
rect 43111 72020 43130 72076
rect 43036 71996 43130 72020
rect 43036 71940 43055 71996
rect 43111 71940 43130 71996
rect 43036 71912 43130 71940
rect 45926 72236 46020 72264
rect 45926 72180 45945 72236
rect 46001 72180 46020 72236
rect 45926 72156 46020 72180
rect 45926 72100 45945 72156
rect 46001 72100 46020 72156
rect 45926 72076 46020 72100
rect 45926 72020 45945 72076
rect 46001 72020 46020 72076
rect 45926 71996 46020 72020
rect 45926 71940 45945 71996
rect 46001 71940 46020 71996
rect 45926 71912 46020 71940
rect 48873 72236 48967 72264
rect 48873 72180 48892 72236
rect 48948 72180 48967 72236
rect 48873 72156 48967 72180
rect 48873 72100 48892 72156
rect 48948 72100 48967 72156
rect 48873 72076 48967 72100
rect 48873 72020 48892 72076
rect 48948 72020 48967 72076
rect 48873 71996 48967 72020
rect 48873 71940 48892 71996
rect 48948 71940 48967 71996
rect 48873 71912 48967 71940
rect 49722 72236 49922 72264
rect 49722 72180 49754 72236
rect 49810 72180 49834 72236
rect 49890 72180 49922 72236
rect 49722 72156 49922 72180
rect 49722 72100 49754 72156
rect 49810 72100 49834 72156
rect 49890 72100 49922 72156
rect 49722 72076 49922 72100
rect 49722 72020 49754 72076
rect 49810 72020 49834 72076
rect 49890 72020 49922 72076
rect 49722 71996 49922 72020
rect 49722 71940 49754 71996
rect 49810 71940 49834 71996
rect 49890 71940 49922 71996
rect 49722 71912 49922 71940
rect 53012 72236 53140 72264
rect 53012 72180 53048 72236
rect 53104 72180 53140 72236
rect 53012 72156 53140 72180
rect 53012 72100 53048 72156
rect 53104 72100 53140 72156
rect 53012 72076 53140 72100
rect 53012 72020 53048 72076
rect 53104 72020 53140 72076
rect 53012 71996 53140 72020
rect 53012 71940 53048 71996
rect 53104 71940 53140 71996
rect 53012 71912 53140 71940
rect 53170 72236 53298 72264
rect 53170 72180 53206 72236
rect 53262 72180 53298 72236
rect 53170 72156 53298 72180
rect 53170 72100 53206 72156
rect 53262 72100 53298 72156
rect 53170 72076 53298 72100
rect 53170 72020 53206 72076
rect 53262 72020 53298 72076
rect 53170 71996 53298 72020
rect 53170 71940 53206 71996
rect 53262 71940 53298 71996
rect 53170 71912 53298 71940
rect 53526 72236 53654 72264
rect 53526 72180 53562 72236
rect 53618 72180 53654 72236
rect 53526 72156 53654 72180
rect 53526 72100 53562 72156
rect 53618 72100 53654 72156
rect 53526 72076 53654 72100
rect 53526 72020 53562 72076
rect 53618 72020 53654 72076
rect 53526 71996 53654 72020
rect 53526 71940 53562 71996
rect 53618 71940 53654 71996
rect 53526 71912 53654 71940
rect 54844 72236 54972 72264
rect 54844 72180 54880 72236
rect 54936 72180 54972 72236
rect 54844 72156 54972 72180
rect 54844 72100 54880 72156
rect 54936 72100 54972 72156
rect 54844 72076 54972 72100
rect 54844 72020 54880 72076
rect 54936 72020 54972 72076
rect 54844 71996 54972 72020
rect 54844 71940 54880 71996
rect 54936 71940 54972 71996
rect 54844 71912 54972 71940
rect 55437 72236 55565 72264
rect 55437 72180 55473 72236
rect 55529 72180 55565 72236
rect 55437 72156 55565 72180
rect 55437 72100 55473 72156
rect 55529 72100 55565 72156
rect 55437 72076 55565 72100
rect 55437 72020 55473 72076
rect 55529 72020 55565 72076
rect 55437 71996 55565 72020
rect 55437 71940 55473 71996
rect 55529 71940 55565 71996
rect 55437 71912 55565 71940
rect 56583 72236 56711 72264
rect 56583 72180 56619 72236
rect 56675 72180 56711 72236
rect 56583 72156 56711 72180
rect 56583 72100 56619 72156
rect 56675 72100 56711 72156
rect 56583 72076 56711 72100
rect 56583 72020 56619 72076
rect 56675 72020 56711 72076
rect 56583 71996 56711 72020
rect 56583 71940 56619 71996
rect 56675 71940 56711 71996
rect 56583 71912 56711 71940
rect 58033 72236 58213 72264
rect 58033 72180 58055 72236
rect 58111 72180 58135 72236
rect 58191 72180 58213 72236
rect 58033 72156 58213 72180
rect 58033 72100 58055 72156
rect 58111 72100 58135 72156
rect 58191 72100 58213 72156
rect 58033 72076 58213 72100
rect 58033 72020 58055 72076
rect 58111 72020 58135 72076
rect 58191 72020 58213 72076
rect 58033 71996 58213 72020
rect 58033 71940 58055 71996
rect 58111 71940 58135 71996
rect 58191 71940 58213 71996
rect 58033 71912 58213 71940
rect 59256 72236 59396 72264
rect 59256 72180 59298 72236
rect 59354 72180 59396 72236
rect 59256 72156 59396 72180
rect 59256 72100 59298 72156
rect 59354 72100 59396 72156
rect 59256 72076 59396 72100
rect 59256 72020 59298 72076
rect 59354 72020 59396 72076
rect 59256 71996 59396 72020
rect 59256 71940 59298 71996
rect 59354 71940 59396 71996
rect 59256 71912 59396 71940
rect 59426 72236 59542 72264
rect 59426 72180 59456 72236
rect 59512 72180 59542 72236
rect 59426 72156 59542 72180
rect 59426 72100 59456 72156
rect 59512 72100 59542 72156
rect 59426 72076 59542 72100
rect 59426 72020 59456 72076
rect 59512 72020 59542 72076
rect 59426 71996 59542 72020
rect 59426 71940 59456 71996
rect 59512 71940 59542 71996
rect 59426 71912 59542 71940
rect 59734 72236 59850 72264
rect 59734 72180 59764 72236
rect 59820 72180 59850 72236
rect 59734 72156 59850 72180
rect 59734 72100 59764 72156
rect 59820 72100 59850 72156
rect 59734 72076 59850 72100
rect 59734 72020 59764 72076
rect 59820 72020 59850 72076
rect 59734 71996 59850 72020
rect 59734 71940 59764 71996
rect 59820 71940 59850 71996
rect 59734 71912 59850 71940
rect 59880 72236 59996 72264
rect 59880 72180 59910 72236
rect 59966 72180 59996 72236
rect 59880 72156 59996 72180
rect 59880 72100 59910 72156
rect 59966 72100 59996 72156
rect 59880 72076 59996 72100
rect 59880 72020 59910 72076
rect 59966 72020 59996 72076
rect 59880 71996 59996 72020
rect 59880 71940 59910 71996
rect 59966 71940 59996 71996
rect 59880 71912 59996 71940
rect 60026 72236 60202 72264
rect 60026 72180 60046 72236
rect 60102 72180 60126 72236
rect 60182 72180 60202 72236
rect 60026 72156 60202 72180
rect 60026 72100 60046 72156
rect 60102 72100 60126 72156
rect 60182 72100 60202 72156
rect 60026 72076 60202 72100
rect 60026 72020 60046 72076
rect 60102 72020 60126 72076
rect 60182 72020 60202 72076
rect 60026 71996 60202 72020
rect 60026 71940 60046 71996
rect 60102 71940 60126 71996
rect 60182 71940 60202 71996
rect 60026 71912 60202 71940
rect 62399 72236 62573 72264
rect 62399 72180 62418 72236
rect 62474 72180 62498 72236
rect 62554 72180 62573 72236
rect 62399 72156 62573 72180
rect 62399 72100 62418 72156
rect 62474 72100 62498 72156
rect 62554 72100 62573 72156
rect 62399 72076 62573 72100
rect 62399 72020 62418 72076
rect 62474 72020 62498 72076
rect 62554 72020 62573 72076
rect 62399 71996 62573 72020
rect 62399 71940 62418 71996
rect 62474 71940 62498 71996
rect 62554 71940 62573 71996
rect 62399 71912 62573 71940
rect 63512 71670 63540 76684
rect 63604 75818 63632 77386
rect 63684 76152 63736 76158
rect 63684 76094 63736 76100
rect 63592 75812 63644 75818
rect 63592 75754 63644 75760
rect 63604 73234 63632 75754
rect 63592 73228 63644 73234
rect 63592 73170 63644 73176
rect 63500 71664 63552 71670
rect 63500 71606 63552 71612
rect 63604 71466 63632 73170
rect 63592 71460 63644 71466
rect 63592 71402 63644 71408
rect 63500 70848 63552 70854
rect 63500 70790 63552 70796
rect 63512 69018 63540 70790
rect 63500 69012 63552 69018
rect 63500 68954 63552 68960
rect 63592 66496 63644 66502
rect 63592 66438 63644 66444
rect 63500 65272 63552 65278
rect 63498 65240 63500 65249
rect 63552 65240 63554 65249
rect 63498 65175 63554 65184
rect 63604 64870 63632 66438
rect 63592 64864 63644 64870
rect 63592 64806 63644 64812
rect 63592 64728 63644 64734
rect 63592 64670 63644 64676
rect 2112 64588 2216 64616
rect 2112 64532 2136 64588
rect 2192 64532 2216 64588
rect 2112 64508 2216 64532
rect 2112 64452 2136 64508
rect 2192 64452 2216 64508
rect 2112 64428 2216 64452
rect 2112 64372 2136 64428
rect 2192 64372 2216 64428
rect 2112 64348 2216 64372
rect 2112 64292 2136 64348
rect 2192 64292 2216 64348
rect 2112 64264 2216 64292
rect 5613 64588 5707 64616
rect 5613 64532 5632 64588
rect 5688 64532 5707 64588
rect 5613 64508 5707 64532
rect 5613 64452 5632 64508
rect 5688 64452 5707 64508
rect 5613 64428 5707 64452
rect 5613 64372 5632 64428
rect 5688 64372 5707 64428
rect 5613 64348 5707 64372
rect 5613 64292 5632 64348
rect 5688 64292 5707 64348
rect 5613 64264 5707 64292
rect 8503 64588 8597 64616
rect 8503 64532 8522 64588
rect 8578 64532 8597 64588
rect 8503 64508 8597 64532
rect 8503 64452 8522 64508
rect 8578 64452 8597 64508
rect 8503 64428 8597 64452
rect 8503 64372 8522 64428
rect 8578 64372 8597 64428
rect 8503 64348 8597 64372
rect 8503 64292 8522 64348
rect 8578 64292 8597 64348
rect 8503 64264 8597 64292
rect 11393 64588 11487 64616
rect 11393 64532 11412 64588
rect 11468 64532 11487 64588
rect 11393 64508 11487 64532
rect 11393 64452 11412 64508
rect 11468 64452 11487 64508
rect 11393 64428 11487 64452
rect 11393 64372 11412 64428
rect 11468 64372 11487 64428
rect 11393 64348 11487 64372
rect 11393 64292 11412 64348
rect 11468 64292 11487 64348
rect 11393 64264 11487 64292
rect 14283 64588 14377 64616
rect 14283 64532 14302 64588
rect 14358 64532 14377 64588
rect 14283 64508 14377 64532
rect 14283 64452 14302 64508
rect 14358 64452 14377 64508
rect 14283 64428 14377 64452
rect 14283 64372 14302 64428
rect 14358 64372 14377 64428
rect 14283 64348 14377 64372
rect 14283 64292 14302 64348
rect 14358 64292 14377 64348
rect 14283 64264 14377 64292
rect 17173 64588 17267 64616
rect 17173 64532 17192 64588
rect 17248 64532 17267 64588
rect 17173 64508 17267 64532
rect 17173 64452 17192 64508
rect 17248 64452 17267 64508
rect 17173 64428 17267 64452
rect 17173 64372 17192 64428
rect 17248 64372 17267 64428
rect 17173 64348 17267 64372
rect 17173 64292 17192 64348
rect 17248 64292 17267 64348
rect 17173 64264 17267 64292
rect 20063 64588 20157 64616
rect 20063 64532 20082 64588
rect 20138 64532 20157 64588
rect 20063 64508 20157 64532
rect 20063 64452 20082 64508
rect 20138 64452 20157 64508
rect 20063 64428 20157 64452
rect 20063 64372 20082 64428
rect 20138 64372 20157 64428
rect 20063 64348 20157 64372
rect 20063 64292 20082 64348
rect 20138 64292 20157 64348
rect 20063 64264 20157 64292
rect 22953 64588 23047 64616
rect 22953 64532 22972 64588
rect 23028 64532 23047 64588
rect 22953 64508 23047 64532
rect 22953 64452 22972 64508
rect 23028 64452 23047 64508
rect 22953 64428 23047 64452
rect 22953 64372 22972 64428
rect 23028 64372 23047 64428
rect 22953 64348 23047 64372
rect 22953 64292 22972 64348
rect 23028 64292 23047 64348
rect 22953 64264 23047 64292
rect 25843 64588 25937 64616
rect 25843 64532 25862 64588
rect 25918 64532 25937 64588
rect 25843 64508 25937 64532
rect 25843 64452 25862 64508
rect 25918 64452 25937 64508
rect 25843 64428 25937 64452
rect 25843 64372 25862 64428
rect 25918 64372 25937 64428
rect 25843 64348 25937 64372
rect 25843 64292 25862 64348
rect 25918 64292 25937 64348
rect 25843 64264 25937 64292
rect 28733 64588 28827 64616
rect 28733 64532 28752 64588
rect 28808 64532 28827 64588
rect 28733 64508 28827 64532
rect 28733 64452 28752 64508
rect 28808 64452 28827 64508
rect 28733 64428 28827 64452
rect 28733 64372 28752 64428
rect 28808 64372 28827 64428
rect 28733 64348 28827 64372
rect 28733 64292 28752 64348
rect 28808 64292 28827 64348
rect 28733 64264 28827 64292
rect 31623 64588 31717 64616
rect 31623 64532 31642 64588
rect 31698 64532 31717 64588
rect 31623 64508 31717 64532
rect 31623 64452 31642 64508
rect 31698 64452 31717 64508
rect 31623 64428 31717 64452
rect 31623 64372 31642 64428
rect 31698 64372 31717 64428
rect 31623 64348 31717 64372
rect 31623 64292 31642 64348
rect 31698 64292 31717 64348
rect 31623 64264 31717 64292
rect 34513 64588 34607 64616
rect 34513 64532 34532 64588
rect 34588 64532 34607 64588
rect 34513 64508 34607 64532
rect 34513 64452 34532 64508
rect 34588 64452 34607 64508
rect 34513 64428 34607 64452
rect 34513 64372 34532 64428
rect 34588 64372 34607 64428
rect 34513 64348 34607 64372
rect 34513 64292 34532 64348
rect 34588 64292 34607 64348
rect 34513 64264 34607 64292
rect 37403 64588 37497 64616
rect 37403 64532 37422 64588
rect 37478 64532 37497 64588
rect 37403 64508 37497 64532
rect 37403 64452 37422 64508
rect 37478 64452 37497 64508
rect 37403 64428 37497 64452
rect 37403 64372 37422 64428
rect 37478 64372 37497 64428
rect 37403 64348 37497 64372
rect 37403 64292 37422 64348
rect 37478 64292 37497 64348
rect 37403 64264 37497 64292
rect 40293 64588 40387 64616
rect 40293 64532 40312 64588
rect 40368 64532 40387 64588
rect 40293 64508 40387 64532
rect 40293 64452 40312 64508
rect 40368 64452 40387 64508
rect 40293 64428 40387 64452
rect 40293 64372 40312 64428
rect 40368 64372 40387 64428
rect 40293 64348 40387 64372
rect 40293 64292 40312 64348
rect 40368 64292 40387 64348
rect 40293 64264 40387 64292
rect 43183 64588 43277 64616
rect 43183 64532 43202 64588
rect 43258 64532 43277 64588
rect 43183 64508 43277 64532
rect 43183 64452 43202 64508
rect 43258 64452 43277 64508
rect 43183 64428 43277 64452
rect 43183 64372 43202 64428
rect 43258 64372 43277 64428
rect 43183 64348 43277 64372
rect 43183 64292 43202 64348
rect 43258 64292 43277 64348
rect 43183 64264 43277 64292
rect 46073 64588 46167 64616
rect 46073 64532 46092 64588
rect 46148 64532 46167 64588
rect 46073 64508 46167 64532
rect 46073 64452 46092 64508
rect 46148 64452 46167 64508
rect 46073 64428 46167 64452
rect 46073 64372 46092 64428
rect 46148 64372 46167 64428
rect 46073 64348 46167 64372
rect 46073 64292 46092 64348
rect 46148 64292 46167 64348
rect 46073 64264 46167 64292
rect 49081 64588 49175 64616
rect 49081 64532 49100 64588
rect 49156 64532 49175 64588
rect 49081 64508 49175 64532
rect 49081 64452 49100 64508
rect 49156 64452 49175 64508
rect 49081 64428 49175 64452
rect 49081 64372 49100 64428
rect 49156 64372 49175 64428
rect 49081 64348 49175 64372
rect 49081 64292 49100 64348
rect 49156 64292 49175 64348
rect 49081 64264 49175 64292
rect 52302 64588 52412 64616
rect 52302 64532 52329 64588
rect 52385 64532 52412 64588
rect 52302 64508 52412 64532
rect 52302 64452 52329 64508
rect 52385 64452 52412 64508
rect 52302 64428 52412 64452
rect 52302 64372 52329 64428
rect 52385 64372 52412 64428
rect 52302 64348 52412 64372
rect 52302 64292 52329 64348
rect 52385 64292 52412 64348
rect 52302 64264 52412 64292
rect 53694 64588 53822 64616
rect 53694 64532 53730 64588
rect 53786 64532 53822 64588
rect 53694 64508 53822 64532
rect 53694 64452 53730 64508
rect 53786 64452 53822 64508
rect 53694 64428 53822 64452
rect 53694 64372 53730 64428
rect 53786 64372 53822 64428
rect 53694 64348 53822 64372
rect 53694 64292 53730 64348
rect 53786 64292 53822 64348
rect 53694 64264 53822 64292
rect 53862 64588 53990 64616
rect 53862 64532 53898 64588
rect 53954 64532 53990 64588
rect 53862 64508 53990 64532
rect 53862 64452 53898 64508
rect 53954 64452 53990 64508
rect 53862 64428 53990 64452
rect 53862 64372 53898 64428
rect 53954 64372 53990 64428
rect 53862 64348 53990 64372
rect 53862 64292 53898 64348
rect 53954 64292 53990 64348
rect 53862 64264 53990 64292
rect 54606 64588 54734 64616
rect 54606 64532 54642 64588
rect 54698 64532 54734 64588
rect 54606 64508 54734 64532
rect 54606 64452 54642 64508
rect 54698 64452 54734 64508
rect 54606 64428 54734 64452
rect 54606 64372 54642 64428
rect 54698 64372 54734 64428
rect 54606 64348 54734 64372
rect 54606 64292 54642 64348
rect 54698 64292 54734 64348
rect 54606 64264 54734 64292
rect 55002 64588 55118 64616
rect 55002 64532 55032 64588
rect 55088 64532 55118 64588
rect 55002 64508 55118 64532
rect 55002 64452 55032 64508
rect 55088 64452 55118 64508
rect 55002 64428 55118 64452
rect 55002 64372 55032 64428
rect 55088 64372 55118 64428
rect 55002 64348 55118 64372
rect 55002 64292 55032 64348
rect 55088 64292 55118 64348
rect 55002 64264 55118 64292
rect 55712 64588 55840 64616
rect 55712 64532 55748 64588
rect 55804 64532 55840 64588
rect 55712 64508 55840 64532
rect 55712 64452 55748 64508
rect 55804 64452 55840 64508
rect 55712 64428 55840 64452
rect 55712 64372 55748 64428
rect 55804 64372 55840 64428
rect 55712 64348 55840 64372
rect 55712 64292 55748 64348
rect 55804 64292 55840 64348
rect 55712 64264 55840 64292
rect 56290 64588 56418 64616
rect 56290 64532 56326 64588
rect 56382 64532 56418 64588
rect 56290 64508 56418 64532
rect 56290 64452 56326 64508
rect 56382 64452 56418 64508
rect 56290 64428 56418 64452
rect 56290 64372 56326 64428
rect 56382 64372 56418 64428
rect 56290 64348 56418 64372
rect 56290 64292 56326 64348
rect 56382 64292 56418 64348
rect 56290 64264 56418 64292
rect 56741 64588 56857 64616
rect 56741 64532 56771 64588
rect 56827 64532 56857 64588
rect 56741 64508 56857 64532
rect 56741 64452 56771 64508
rect 56827 64452 56857 64508
rect 56741 64428 56857 64452
rect 56741 64372 56771 64428
rect 56827 64372 56857 64428
rect 56741 64348 56857 64372
rect 56741 64292 56771 64348
rect 56827 64292 56857 64348
rect 56741 64264 56857 64292
rect 57045 64588 57161 64616
rect 57045 64532 57075 64588
rect 57131 64532 57161 64588
rect 57045 64508 57161 64532
rect 57045 64452 57075 64508
rect 57131 64452 57161 64508
rect 57045 64428 57161 64452
rect 57045 64372 57075 64428
rect 57131 64372 57161 64428
rect 57045 64348 57161 64372
rect 57045 64292 57075 64348
rect 57131 64292 57161 64348
rect 57045 64264 57161 64292
rect 57887 64588 58003 64616
rect 57887 64532 57917 64588
rect 57973 64532 58003 64588
rect 57887 64508 58003 64532
rect 57887 64452 57917 64508
rect 57973 64452 58003 64508
rect 57887 64428 58003 64452
rect 57887 64372 57917 64428
rect 57973 64372 58003 64428
rect 57887 64348 58003 64372
rect 57887 64292 57917 64348
rect 57973 64292 58003 64348
rect 57887 64264 58003 64292
rect 58553 64588 58617 64616
rect 58553 64532 58557 64588
rect 58613 64532 58617 64588
rect 58553 64508 58617 64532
rect 58553 64452 58557 64508
rect 58613 64452 58617 64508
rect 58553 64428 58617 64452
rect 58553 64372 58557 64428
rect 58613 64372 58617 64428
rect 58553 64348 58617 64372
rect 58553 64292 58557 64348
rect 58613 64292 58617 64348
rect 58553 64264 58617 64292
rect 59110 64588 59226 64616
rect 59110 64532 59140 64588
rect 59196 64532 59226 64588
rect 59110 64508 59226 64532
rect 59110 64452 59140 64508
rect 59196 64452 59226 64508
rect 59110 64428 59226 64452
rect 59110 64372 59140 64428
rect 59196 64372 59226 64428
rect 59110 64348 59226 64372
rect 59110 64292 59140 64348
rect 59196 64292 59226 64348
rect 59110 64264 59226 64292
rect 60388 64588 60504 64616
rect 60388 64532 60418 64588
rect 60474 64532 60504 64588
rect 60388 64508 60504 64532
rect 60388 64452 60418 64508
rect 60474 64452 60504 64508
rect 60388 64428 60504 64452
rect 60388 64372 60418 64428
rect 60474 64372 60504 64428
rect 60388 64348 60504 64372
rect 60388 64292 60418 64348
rect 60474 64292 60504 64348
rect 60388 64264 60504 64292
rect 60546 64588 60662 64616
rect 60546 64532 60576 64588
rect 60632 64532 60662 64588
rect 60546 64508 60662 64532
rect 60546 64452 60576 64508
rect 60632 64452 60662 64508
rect 60546 64428 60662 64452
rect 60546 64372 60576 64428
rect 60632 64372 60662 64428
rect 60546 64348 60662 64372
rect 60546 64292 60576 64348
rect 60632 64292 60662 64348
rect 60546 64264 60662 64292
rect 62601 64588 62775 64616
rect 62601 64532 62620 64588
rect 62676 64532 62700 64588
rect 62756 64532 62775 64588
rect 62601 64508 62775 64532
rect 62601 64452 62620 64508
rect 62676 64452 62700 64508
rect 62756 64452 62775 64508
rect 62601 64428 62775 64452
rect 62601 64372 62620 64428
rect 62676 64372 62700 64428
rect 62756 64372 62775 64428
rect 62601 64348 62775 64372
rect 62601 64292 62620 64348
rect 62676 64292 62700 64348
rect 62756 64292 62775 64348
rect 62601 64264 62775 64292
rect 63500 63232 63552 63238
rect 63498 63200 63500 63209
rect 63552 63200 63554 63209
rect 63498 63135 63554 63144
rect 2244 62236 2444 62264
rect 2244 62180 2276 62236
rect 2332 62180 2356 62236
rect 2412 62180 2444 62236
rect 2244 62156 2444 62180
rect 2244 62100 2276 62156
rect 2332 62100 2356 62156
rect 2412 62100 2444 62156
rect 2244 62076 2444 62100
rect 2244 62020 2276 62076
rect 2332 62020 2356 62076
rect 2412 62020 2444 62076
rect 2244 61996 2444 62020
rect 2244 61940 2276 61996
rect 2332 61940 2356 61996
rect 2412 61940 2444 61996
rect 2244 61912 2444 61940
rect 5466 62236 5560 62264
rect 5466 62180 5485 62236
rect 5541 62180 5560 62236
rect 5466 62156 5560 62180
rect 5466 62100 5485 62156
rect 5541 62100 5560 62156
rect 5466 62076 5560 62100
rect 5466 62020 5485 62076
rect 5541 62020 5560 62076
rect 5466 61996 5560 62020
rect 5466 61940 5485 61996
rect 5541 61940 5560 61996
rect 5466 61912 5560 61940
rect 8356 62236 8450 62264
rect 8356 62180 8375 62236
rect 8431 62180 8450 62236
rect 8356 62156 8450 62180
rect 8356 62100 8375 62156
rect 8431 62100 8450 62156
rect 8356 62076 8450 62100
rect 8356 62020 8375 62076
rect 8431 62020 8450 62076
rect 8356 61996 8450 62020
rect 8356 61940 8375 61996
rect 8431 61940 8450 61996
rect 8356 61912 8450 61940
rect 11246 62236 11340 62264
rect 11246 62180 11265 62236
rect 11321 62180 11340 62236
rect 11246 62156 11340 62180
rect 11246 62100 11265 62156
rect 11321 62100 11340 62156
rect 11246 62076 11340 62100
rect 11246 62020 11265 62076
rect 11321 62020 11340 62076
rect 11246 61996 11340 62020
rect 11246 61940 11265 61996
rect 11321 61940 11340 61996
rect 11246 61912 11340 61940
rect 14136 62236 14230 62264
rect 14136 62180 14155 62236
rect 14211 62180 14230 62236
rect 14136 62156 14230 62180
rect 14136 62100 14155 62156
rect 14211 62100 14230 62156
rect 14136 62076 14230 62100
rect 14136 62020 14155 62076
rect 14211 62020 14230 62076
rect 14136 61996 14230 62020
rect 14136 61940 14155 61996
rect 14211 61940 14230 61996
rect 14136 61912 14230 61940
rect 17026 62236 17120 62264
rect 17026 62180 17045 62236
rect 17101 62180 17120 62236
rect 17026 62156 17120 62180
rect 17026 62100 17045 62156
rect 17101 62100 17120 62156
rect 17026 62076 17120 62100
rect 17026 62020 17045 62076
rect 17101 62020 17120 62076
rect 17026 61996 17120 62020
rect 17026 61940 17045 61996
rect 17101 61940 17120 61996
rect 17026 61912 17120 61940
rect 19916 62236 20010 62264
rect 19916 62180 19935 62236
rect 19991 62180 20010 62236
rect 19916 62156 20010 62180
rect 19916 62100 19935 62156
rect 19991 62100 20010 62156
rect 19916 62076 20010 62100
rect 19916 62020 19935 62076
rect 19991 62020 20010 62076
rect 19916 61996 20010 62020
rect 19916 61940 19935 61996
rect 19991 61940 20010 61996
rect 19916 61912 20010 61940
rect 22806 62236 22900 62264
rect 22806 62180 22825 62236
rect 22881 62180 22900 62236
rect 22806 62156 22900 62180
rect 22806 62100 22825 62156
rect 22881 62100 22900 62156
rect 22806 62076 22900 62100
rect 22806 62020 22825 62076
rect 22881 62020 22900 62076
rect 22806 61996 22900 62020
rect 22806 61940 22825 61996
rect 22881 61940 22900 61996
rect 22806 61912 22900 61940
rect 25696 62236 25790 62264
rect 25696 62180 25715 62236
rect 25771 62180 25790 62236
rect 25696 62156 25790 62180
rect 25696 62100 25715 62156
rect 25771 62100 25790 62156
rect 25696 62076 25790 62100
rect 25696 62020 25715 62076
rect 25771 62020 25790 62076
rect 25696 61996 25790 62020
rect 25696 61940 25715 61996
rect 25771 61940 25790 61996
rect 25696 61912 25790 61940
rect 28586 62236 28680 62264
rect 28586 62180 28605 62236
rect 28661 62180 28680 62236
rect 28586 62156 28680 62180
rect 28586 62100 28605 62156
rect 28661 62100 28680 62156
rect 28586 62076 28680 62100
rect 28586 62020 28605 62076
rect 28661 62020 28680 62076
rect 28586 61996 28680 62020
rect 28586 61940 28605 61996
rect 28661 61940 28680 61996
rect 28586 61912 28680 61940
rect 31476 62236 31570 62264
rect 31476 62180 31495 62236
rect 31551 62180 31570 62236
rect 31476 62156 31570 62180
rect 31476 62100 31495 62156
rect 31551 62100 31570 62156
rect 31476 62076 31570 62100
rect 31476 62020 31495 62076
rect 31551 62020 31570 62076
rect 31476 61996 31570 62020
rect 31476 61940 31495 61996
rect 31551 61940 31570 61996
rect 31476 61912 31570 61940
rect 34366 62236 34460 62264
rect 34366 62180 34385 62236
rect 34441 62180 34460 62236
rect 34366 62156 34460 62180
rect 34366 62100 34385 62156
rect 34441 62100 34460 62156
rect 34366 62076 34460 62100
rect 34366 62020 34385 62076
rect 34441 62020 34460 62076
rect 34366 61996 34460 62020
rect 34366 61940 34385 61996
rect 34441 61940 34460 61996
rect 34366 61912 34460 61940
rect 37256 62236 37350 62264
rect 37256 62180 37275 62236
rect 37331 62180 37350 62236
rect 37256 62156 37350 62180
rect 37256 62100 37275 62156
rect 37331 62100 37350 62156
rect 37256 62076 37350 62100
rect 37256 62020 37275 62076
rect 37331 62020 37350 62076
rect 37256 61996 37350 62020
rect 37256 61940 37275 61996
rect 37331 61940 37350 61996
rect 37256 61912 37350 61940
rect 40146 62236 40240 62264
rect 40146 62180 40165 62236
rect 40221 62180 40240 62236
rect 40146 62156 40240 62180
rect 40146 62100 40165 62156
rect 40221 62100 40240 62156
rect 40146 62076 40240 62100
rect 40146 62020 40165 62076
rect 40221 62020 40240 62076
rect 40146 61996 40240 62020
rect 40146 61940 40165 61996
rect 40221 61940 40240 61996
rect 40146 61912 40240 61940
rect 43036 62236 43130 62264
rect 43036 62180 43055 62236
rect 43111 62180 43130 62236
rect 43036 62156 43130 62180
rect 43036 62100 43055 62156
rect 43111 62100 43130 62156
rect 43036 62076 43130 62100
rect 43036 62020 43055 62076
rect 43111 62020 43130 62076
rect 43036 61996 43130 62020
rect 43036 61940 43055 61996
rect 43111 61940 43130 61996
rect 43036 61912 43130 61940
rect 45926 62236 46020 62264
rect 45926 62180 45945 62236
rect 46001 62180 46020 62236
rect 45926 62156 46020 62180
rect 45926 62100 45945 62156
rect 46001 62100 46020 62156
rect 45926 62076 46020 62100
rect 45926 62020 45945 62076
rect 46001 62020 46020 62076
rect 45926 61996 46020 62020
rect 45926 61940 45945 61996
rect 46001 61940 46020 61996
rect 45926 61912 46020 61940
rect 48873 62236 48967 62264
rect 48873 62180 48892 62236
rect 48948 62180 48967 62236
rect 48873 62156 48967 62180
rect 48873 62100 48892 62156
rect 48948 62100 48967 62156
rect 48873 62076 48967 62100
rect 48873 62020 48892 62076
rect 48948 62020 48967 62076
rect 48873 61996 48967 62020
rect 48873 61940 48892 61996
rect 48948 61940 48967 61996
rect 48873 61912 48967 61940
rect 49722 62236 49922 62264
rect 49722 62180 49754 62236
rect 49810 62180 49834 62236
rect 49890 62180 49922 62236
rect 49722 62156 49922 62180
rect 49722 62100 49754 62156
rect 49810 62100 49834 62156
rect 49890 62100 49922 62156
rect 49722 62076 49922 62100
rect 49722 62020 49754 62076
rect 49810 62020 49834 62076
rect 49890 62020 49922 62076
rect 49722 61996 49922 62020
rect 49722 61940 49754 61996
rect 49810 61940 49834 61996
rect 49890 61940 49922 61996
rect 49722 61912 49922 61940
rect 53012 62236 53140 62264
rect 53012 62180 53048 62236
rect 53104 62180 53140 62236
rect 53012 62156 53140 62180
rect 53012 62100 53048 62156
rect 53104 62100 53140 62156
rect 53012 62076 53140 62100
rect 53012 62020 53048 62076
rect 53104 62020 53140 62076
rect 53012 61996 53140 62020
rect 53012 61940 53048 61996
rect 53104 61940 53140 61996
rect 53012 61912 53140 61940
rect 53170 62236 53298 62264
rect 53170 62180 53206 62236
rect 53262 62180 53298 62236
rect 53170 62156 53298 62180
rect 53170 62100 53206 62156
rect 53262 62100 53298 62156
rect 53170 62076 53298 62100
rect 53170 62020 53206 62076
rect 53262 62020 53298 62076
rect 53170 61996 53298 62020
rect 53170 61940 53206 61996
rect 53262 61940 53298 61996
rect 53170 61912 53298 61940
rect 53526 62236 53654 62264
rect 53526 62180 53562 62236
rect 53618 62180 53654 62236
rect 53526 62156 53654 62180
rect 53526 62100 53562 62156
rect 53618 62100 53654 62156
rect 53526 62076 53654 62100
rect 53526 62020 53562 62076
rect 53618 62020 53654 62076
rect 53526 61996 53654 62020
rect 53526 61940 53562 61996
rect 53618 61940 53654 61996
rect 53526 61912 53654 61940
rect 54844 62236 54972 62264
rect 54844 62180 54880 62236
rect 54936 62180 54972 62236
rect 54844 62156 54972 62180
rect 54844 62100 54880 62156
rect 54936 62100 54972 62156
rect 54844 62076 54972 62100
rect 54844 62020 54880 62076
rect 54936 62020 54972 62076
rect 54844 61996 54972 62020
rect 54844 61940 54880 61996
rect 54936 61940 54972 61996
rect 54844 61912 54972 61940
rect 55437 62236 55565 62264
rect 55437 62180 55473 62236
rect 55529 62180 55565 62236
rect 55437 62156 55565 62180
rect 55437 62100 55473 62156
rect 55529 62100 55565 62156
rect 55437 62076 55565 62100
rect 55437 62020 55473 62076
rect 55529 62020 55565 62076
rect 55437 61996 55565 62020
rect 55437 61940 55473 61996
rect 55529 61940 55565 61996
rect 55437 61912 55565 61940
rect 56583 62236 56711 62264
rect 56583 62180 56619 62236
rect 56675 62180 56711 62236
rect 56583 62156 56711 62180
rect 56583 62100 56619 62156
rect 56675 62100 56711 62156
rect 56583 62076 56711 62100
rect 56583 62020 56619 62076
rect 56675 62020 56711 62076
rect 56583 61996 56711 62020
rect 56583 61940 56619 61996
rect 56675 61940 56711 61996
rect 56583 61912 56711 61940
rect 58033 62236 58213 62264
rect 58033 62180 58055 62236
rect 58111 62180 58135 62236
rect 58191 62180 58213 62236
rect 58033 62156 58213 62180
rect 58033 62100 58055 62156
rect 58111 62100 58135 62156
rect 58191 62100 58213 62156
rect 58033 62076 58213 62100
rect 58033 62020 58055 62076
rect 58111 62020 58135 62076
rect 58191 62020 58213 62076
rect 58033 61996 58213 62020
rect 58033 61940 58055 61996
rect 58111 61940 58135 61996
rect 58191 61940 58213 61996
rect 58033 61912 58213 61940
rect 59256 62236 59396 62264
rect 59256 62180 59298 62236
rect 59354 62180 59396 62236
rect 59256 62156 59396 62180
rect 59256 62100 59298 62156
rect 59354 62100 59396 62156
rect 59256 62076 59396 62100
rect 59256 62020 59298 62076
rect 59354 62020 59396 62076
rect 59256 61996 59396 62020
rect 59256 61940 59298 61996
rect 59354 61940 59396 61996
rect 59256 61912 59396 61940
rect 59426 62236 59542 62264
rect 59426 62180 59456 62236
rect 59512 62180 59542 62236
rect 59426 62156 59542 62180
rect 59426 62100 59456 62156
rect 59512 62100 59542 62156
rect 59426 62076 59542 62100
rect 59426 62020 59456 62076
rect 59512 62020 59542 62076
rect 59426 61996 59542 62020
rect 59426 61940 59456 61996
rect 59512 61940 59542 61996
rect 59426 61912 59542 61940
rect 59734 62236 59850 62264
rect 59734 62180 59764 62236
rect 59820 62180 59850 62236
rect 59734 62156 59850 62180
rect 59734 62100 59764 62156
rect 59820 62100 59850 62156
rect 59734 62076 59850 62100
rect 59734 62020 59764 62076
rect 59820 62020 59850 62076
rect 59734 61996 59850 62020
rect 59734 61940 59764 61996
rect 59820 61940 59850 61996
rect 59734 61912 59850 61940
rect 59880 62236 59996 62264
rect 59880 62180 59910 62236
rect 59966 62180 59996 62236
rect 59880 62156 59996 62180
rect 59880 62100 59910 62156
rect 59966 62100 59996 62156
rect 59880 62076 59996 62100
rect 59880 62020 59910 62076
rect 59966 62020 59996 62076
rect 59880 61996 59996 62020
rect 59880 61940 59910 61996
rect 59966 61940 59996 61996
rect 59880 61912 59996 61940
rect 60026 62236 60202 62264
rect 60026 62180 60046 62236
rect 60102 62180 60126 62236
rect 60182 62180 60202 62236
rect 60026 62156 60202 62180
rect 60026 62100 60046 62156
rect 60102 62100 60126 62156
rect 60182 62100 60202 62156
rect 60026 62076 60202 62100
rect 60026 62020 60046 62076
rect 60102 62020 60126 62076
rect 60182 62020 60202 62076
rect 60026 61996 60202 62020
rect 60026 61940 60046 61996
rect 60102 61940 60126 61996
rect 60182 61940 60202 61996
rect 60026 61912 60202 61940
rect 62399 62236 62573 62264
rect 62399 62180 62418 62236
rect 62474 62180 62498 62236
rect 62554 62180 62573 62236
rect 62399 62156 62573 62180
rect 62399 62100 62418 62156
rect 62474 62100 62498 62156
rect 62554 62100 62573 62156
rect 62399 62076 62573 62100
rect 62399 62020 62418 62076
rect 62474 62020 62498 62076
rect 62554 62020 62573 62076
rect 62399 61996 62573 62020
rect 62399 61940 62418 61996
rect 62474 61940 62498 61996
rect 62554 61940 62573 61996
rect 62399 61912 62573 61940
rect 63500 61056 63552 61062
rect 63498 61024 63500 61033
rect 63552 61024 63554 61033
rect 63498 60959 63554 60968
rect 63500 58744 63552 58750
rect 63498 58712 63500 58721
rect 63552 58712 63554 58721
rect 63498 58647 63554 58656
rect 63500 56704 63552 56710
rect 63498 56672 63500 56681
rect 63552 56672 63554 56681
rect 63498 56607 63554 56616
rect 63498 54768 63554 54777
rect 63498 54703 63554 54712
rect 63512 54670 63540 54703
rect 63500 54664 63552 54670
rect 2112 54588 2216 54616
rect 2112 54532 2136 54588
rect 2192 54532 2216 54588
rect 2112 54508 2216 54532
rect 2112 54452 2136 54508
rect 2192 54452 2216 54508
rect 2112 54428 2216 54452
rect 2112 54372 2136 54428
rect 2192 54372 2216 54428
rect 2112 54348 2216 54372
rect 2112 54292 2136 54348
rect 2192 54292 2216 54348
rect 2112 54264 2216 54292
rect 5613 54588 5707 54616
rect 5613 54532 5632 54588
rect 5688 54532 5707 54588
rect 5613 54508 5707 54532
rect 5613 54452 5632 54508
rect 5688 54452 5707 54508
rect 5613 54428 5707 54452
rect 5613 54372 5632 54428
rect 5688 54372 5707 54428
rect 5613 54348 5707 54372
rect 5613 54292 5632 54348
rect 5688 54292 5707 54348
rect 5613 54264 5707 54292
rect 8503 54588 8597 54616
rect 8503 54532 8522 54588
rect 8578 54532 8597 54588
rect 8503 54508 8597 54532
rect 8503 54452 8522 54508
rect 8578 54452 8597 54508
rect 8503 54428 8597 54452
rect 8503 54372 8522 54428
rect 8578 54372 8597 54428
rect 8503 54348 8597 54372
rect 8503 54292 8522 54348
rect 8578 54292 8597 54348
rect 8503 54264 8597 54292
rect 11393 54588 11487 54616
rect 11393 54532 11412 54588
rect 11468 54532 11487 54588
rect 11393 54508 11487 54532
rect 11393 54452 11412 54508
rect 11468 54452 11487 54508
rect 11393 54428 11487 54452
rect 11393 54372 11412 54428
rect 11468 54372 11487 54428
rect 11393 54348 11487 54372
rect 11393 54292 11412 54348
rect 11468 54292 11487 54348
rect 11393 54264 11487 54292
rect 14283 54588 14377 54616
rect 14283 54532 14302 54588
rect 14358 54532 14377 54588
rect 14283 54508 14377 54532
rect 14283 54452 14302 54508
rect 14358 54452 14377 54508
rect 14283 54428 14377 54452
rect 14283 54372 14302 54428
rect 14358 54372 14377 54428
rect 14283 54348 14377 54372
rect 14283 54292 14302 54348
rect 14358 54292 14377 54348
rect 14283 54264 14377 54292
rect 17173 54588 17267 54616
rect 17173 54532 17192 54588
rect 17248 54532 17267 54588
rect 17173 54508 17267 54532
rect 17173 54452 17192 54508
rect 17248 54452 17267 54508
rect 17173 54428 17267 54452
rect 17173 54372 17192 54428
rect 17248 54372 17267 54428
rect 17173 54348 17267 54372
rect 17173 54292 17192 54348
rect 17248 54292 17267 54348
rect 17173 54264 17267 54292
rect 20063 54588 20157 54616
rect 20063 54532 20082 54588
rect 20138 54532 20157 54588
rect 20063 54508 20157 54532
rect 20063 54452 20082 54508
rect 20138 54452 20157 54508
rect 20063 54428 20157 54452
rect 20063 54372 20082 54428
rect 20138 54372 20157 54428
rect 20063 54348 20157 54372
rect 20063 54292 20082 54348
rect 20138 54292 20157 54348
rect 20063 54264 20157 54292
rect 22953 54588 23047 54616
rect 22953 54532 22972 54588
rect 23028 54532 23047 54588
rect 22953 54508 23047 54532
rect 22953 54452 22972 54508
rect 23028 54452 23047 54508
rect 22953 54428 23047 54452
rect 22953 54372 22972 54428
rect 23028 54372 23047 54428
rect 22953 54348 23047 54372
rect 22953 54292 22972 54348
rect 23028 54292 23047 54348
rect 22953 54264 23047 54292
rect 25843 54588 25937 54616
rect 25843 54532 25862 54588
rect 25918 54532 25937 54588
rect 25843 54508 25937 54532
rect 25843 54452 25862 54508
rect 25918 54452 25937 54508
rect 25843 54428 25937 54452
rect 25843 54372 25862 54428
rect 25918 54372 25937 54428
rect 25843 54348 25937 54372
rect 25843 54292 25862 54348
rect 25918 54292 25937 54348
rect 25843 54264 25937 54292
rect 28733 54588 28827 54616
rect 28733 54532 28752 54588
rect 28808 54532 28827 54588
rect 28733 54508 28827 54532
rect 28733 54452 28752 54508
rect 28808 54452 28827 54508
rect 28733 54428 28827 54452
rect 28733 54372 28752 54428
rect 28808 54372 28827 54428
rect 28733 54348 28827 54372
rect 28733 54292 28752 54348
rect 28808 54292 28827 54348
rect 28733 54264 28827 54292
rect 31623 54588 31717 54616
rect 31623 54532 31642 54588
rect 31698 54532 31717 54588
rect 31623 54508 31717 54532
rect 31623 54452 31642 54508
rect 31698 54452 31717 54508
rect 31623 54428 31717 54452
rect 31623 54372 31642 54428
rect 31698 54372 31717 54428
rect 31623 54348 31717 54372
rect 31623 54292 31642 54348
rect 31698 54292 31717 54348
rect 31623 54264 31717 54292
rect 34513 54588 34607 54616
rect 34513 54532 34532 54588
rect 34588 54532 34607 54588
rect 34513 54508 34607 54532
rect 34513 54452 34532 54508
rect 34588 54452 34607 54508
rect 34513 54428 34607 54452
rect 34513 54372 34532 54428
rect 34588 54372 34607 54428
rect 34513 54348 34607 54372
rect 34513 54292 34532 54348
rect 34588 54292 34607 54348
rect 34513 54264 34607 54292
rect 37403 54588 37497 54616
rect 37403 54532 37422 54588
rect 37478 54532 37497 54588
rect 37403 54508 37497 54532
rect 37403 54452 37422 54508
rect 37478 54452 37497 54508
rect 37403 54428 37497 54452
rect 37403 54372 37422 54428
rect 37478 54372 37497 54428
rect 37403 54348 37497 54372
rect 37403 54292 37422 54348
rect 37478 54292 37497 54348
rect 37403 54264 37497 54292
rect 40293 54588 40387 54616
rect 40293 54532 40312 54588
rect 40368 54532 40387 54588
rect 40293 54508 40387 54532
rect 40293 54452 40312 54508
rect 40368 54452 40387 54508
rect 40293 54428 40387 54452
rect 40293 54372 40312 54428
rect 40368 54372 40387 54428
rect 40293 54348 40387 54372
rect 40293 54292 40312 54348
rect 40368 54292 40387 54348
rect 40293 54264 40387 54292
rect 43183 54588 43277 54616
rect 43183 54532 43202 54588
rect 43258 54532 43277 54588
rect 43183 54508 43277 54532
rect 43183 54452 43202 54508
rect 43258 54452 43277 54508
rect 43183 54428 43277 54452
rect 43183 54372 43202 54428
rect 43258 54372 43277 54428
rect 43183 54348 43277 54372
rect 43183 54292 43202 54348
rect 43258 54292 43277 54348
rect 43183 54264 43277 54292
rect 46073 54588 46167 54616
rect 46073 54532 46092 54588
rect 46148 54532 46167 54588
rect 46073 54508 46167 54532
rect 46073 54452 46092 54508
rect 46148 54452 46167 54508
rect 46073 54428 46167 54452
rect 46073 54372 46092 54428
rect 46148 54372 46167 54428
rect 46073 54348 46167 54372
rect 46073 54292 46092 54348
rect 46148 54292 46167 54348
rect 46073 54264 46167 54292
rect 49081 54588 49175 54616
rect 49081 54532 49100 54588
rect 49156 54532 49175 54588
rect 49081 54508 49175 54532
rect 49081 54452 49100 54508
rect 49156 54452 49175 54508
rect 49081 54428 49175 54452
rect 49081 54372 49100 54428
rect 49156 54372 49175 54428
rect 49081 54348 49175 54372
rect 49081 54292 49100 54348
rect 49156 54292 49175 54348
rect 49081 54264 49175 54292
rect 52302 54588 52412 54616
rect 52302 54532 52329 54588
rect 52385 54532 52412 54588
rect 52302 54508 52412 54532
rect 52302 54452 52329 54508
rect 52385 54452 52412 54508
rect 52302 54428 52412 54452
rect 52302 54372 52329 54428
rect 52385 54372 52412 54428
rect 52302 54348 52412 54372
rect 52302 54292 52329 54348
rect 52385 54292 52412 54348
rect 52302 54264 52412 54292
rect 53694 54588 53822 54616
rect 53694 54532 53730 54588
rect 53786 54532 53822 54588
rect 53694 54508 53822 54532
rect 53694 54452 53730 54508
rect 53786 54452 53822 54508
rect 53694 54428 53822 54452
rect 53694 54372 53730 54428
rect 53786 54372 53822 54428
rect 53694 54348 53822 54372
rect 53694 54292 53730 54348
rect 53786 54292 53822 54348
rect 53694 54264 53822 54292
rect 53862 54588 53990 54616
rect 53862 54532 53898 54588
rect 53954 54532 53990 54588
rect 53862 54508 53990 54532
rect 53862 54452 53898 54508
rect 53954 54452 53990 54508
rect 53862 54428 53990 54452
rect 53862 54372 53898 54428
rect 53954 54372 53990 54428
rect 53862 54348 53990 54372
rect 53862 54292 53898 54348
rect 53954 54292 53990 54348
rect 53862 54264 53990 54292
rect 54606 54588 54734 54616
rect 54606 54532 54642 54588
rect 54698 54532 54734 54588
rect 54606 54508 54734 54532
rect 54606 54452 54642 54508
rect 54698 54452 54734 54508
rect 54606 54428 54734 54452
rect 54606 54372 54642 54428
rect 54698 54372 54734 54428
rect 54606 54348 54734 54372
rect 54606 54292 54642 54348
rect 54698 54292 54734 54348
rect 54606 54264 54734 54292
rect 55002 54588 55118 54616
rect 55002 54532 55032 54588
rect 55088 54532 55118 54588
rect 55002 54508 55118 54532
rect 55002 54452 55032 54508
rect 55088 54452 55118 54508
rect 55002 54428 55118 54452
rect 55002 54372 55032 54428
rect 55088 54372 55118 54428
rect 55002 54348 55118 54372
rect 55002 54292 55032 54348
rect 55088 54292 55118 54348
rect 55002 54264 55118 54292
rect 55712 54588 55840 54616
rect 55712 54532 55748 54588
rect 55804 54532 55840 54588
rect 55712 54508 55840 54532
rect 55712 54452 55748 54508
rect 55804 54452 55840 54508
rect 55712 54428 55840 54452
rect 55712 54372 55748 54428
rect 55804 54372 55840 54428
rect 55712 54348 55840 54372
rect 55712 54292 55748 54348
rect 55804 54292 55840 54348
rect 55712 54264 55840 54292
rect 56290 54588 56418 54616
rect 56290 54532 56326 54588
rect 56382 54532 56418 54588
rect 56290 54508 56418 54532
rect 56290 54452 56326 54508
rect 56382 54452 56418 54508
rect 56290 54428 56418 54452
rect 56290 54372 56326 54428
rect 56382 54372 56418 54428
rect 56290 54348 56418 54372
rect 56290 54292 56326 54348
rect 56382 54292 56418 54348
rect 56290 54264 56418 54292
rect 56741 54588 56857 54616
rect 56741 54532 56771 54588
rect 56827 54532 56857 54588
rect 56741 54508 56857 54532
rect 56741 54452 56771 54508
rect 56827 54452 56857 54508
rect 56741 54428 56857 54452
rect 56741 54372 56771 54428
rect 56827 54372 56857 54428
rect 56741 54348 56857 54372
rect 56741 54292 56771 54348
rect 56827 54292 56857 54348
rect 56741 54264 56857 54292
rect 57045 54588 57161 54616
rect 57045 54532 57075 54588
rect 57131 54532 57161 54588
rect 57045 54508 57161 54532
rect 57045 54452 57075 54508
rect 57131 54452 57161 54508
rect 57045 54428 57161 54452
rect 57045 54372 57075 54428
rect 57131 54372 57161 54428
rect 57045 54348 57161 54372
rect 57045 54292 57075 54348
rect 57131 54292 57161 54348
rect 57045 54264 57161 54292
rect 57887 54588 58003 54616
rect 57887 54532 57917 54588
rect 57973 54532 58003 54588
rect 57887 54508 58003 54532
rect 57887 54452 57917 54508
rect 57973 54452 58003 54508
rect 57887 54428 58003 54452
rect 57887 54372 57917 54428
rect 57973 54372 58003 54428
rect 57887 54348 58003 54372
rect 57887 54292 57917 54348
rect 57973 54292 58003 54348
rect 57887 54264 58003 54292
rect 58553 54588 58617 54616
rect 58553 54532 58557 54588
rect 58613 54532 58617 54588
rect 58553 54508 58617 54532
rect 58553 54452 58557 54508
rect 58613 54452 58617 54508
rect 58553 54428 58617 54452
rect 58553 54372 58557 54428
rect 58613 54372 58617 54428
rect 58553 54348 58617 54372
rect 58553 54292 58557 54348
rect 58613 54292 58617 54348
rect 58553 54264 58617 54292
rect 59110 54588 59226 54616
rect 59110 54532 59140 54588
rect 59196 54532 59226 54588
rect 59110 54508 59226 54532
rect 59110 54452 59140 54508
rect 59196 54452 59226 54508
rect 59110 54428 59226 54452
rect 59110 54372 59140 54428
rect 59196 54372 59226 54428
rect 59110 54348 59226 54372
rect 59110 54292 59140 54348
rect 59196 54292 59226 54348
rect 59110 54264 59226 54292
rect 60388 54588 60504 54616
rect 60388 54532 60418 54588
rect 60474 54532 60504 54588
rect 60388 54508 60504 54532
rect 60388 54452 60418 54508
rect 60474 54452 60504 54508
rect 60388 54428 60504 54452
rect 60388 54372 60418 54428
rect 60474 54372 60504 54428
rect 60388 54348 60504 54372
rect 60388 54292 60418 54348
rect 60474 54292 60504 54348
rect 60388 54264 60504 54292
rect 60546 54588 60662 54616
rect 60546 54532 60576 54588
rect 60632 54532 60662 54588
rect 60546 54508 60662 54532
rect 60546 54452 60576 54508
rect 60632 54452 60662 54508
rect 60546 54428 60662 54452
rect 60546 54372 60576 54428
rect 60632 54372 60662 54428
rect 60546 54348 60662 54372
rect 60546 54292 60576 54348
rect 60632 54292 60662 54348
rect 60546 54264 60662 54292
rect 62601 54588 62775 54616
rect 63500 54606 63552 54612
rect 62601 54532 62620 54588
rect 62676 54532 62700 54588
rect 62756 54532 62775 54588
rect 62601 54508 62775 54532
rect 62601 54452 62620 54508
rect 62676 54452 62700 54508
rect 62756 54452 62775 54508
rect 62601 54428 62775 54452
rect 62601 54372 62620 54428
rect 62676 54372 62700 54428
rect 62756 54372 62775 54428
rect 62601 54348 62775 54372
rect 62601 54292 62620 54348
rect 62676 54292 62700 54348
rect 62756 54292 62775 54348
rect 62601 54264 62775 54292
rect 63500 52624 63552 52630
rect 63500 52566 63552 52572
rect 2244 52236 2444 52264
rect 2244 52180 2276 52236
rect 2332 52180 2356 52236
rect 2412 52180 2444 52236
rect 2244 52156 2444 52180
rect 2244 52100 2276 52156
rect 2332 52100 2356 52156
rect 2412 52100 2444 52156
rect 2244 52076 2444 52100
rect 2244 52020 2276 52076
rect 2332 52020 2356 52076
rect 2412 52020 2444 52076
rect 2244 51996 2444 52020
rect 2244 51940 2276 51996
rect 2332 51940 2356 51996
rect 2412 51940 2444 51996
rect 2244 51912 2444 51940
rect 5466 52236 5560 52264
rect 5466 52180 5485 52236
rect 5541 52180 5560 52236
rect 5466 52156 5560 52180
rect 5466 52100 5485 52156
rect 5541 52100 5560 52156
rect 5466 52076 5560 52100
rect 5466 52020 5485 52076
rect 5541 52020 5560 52076
rect 5466 51996 5560 52020
rect 5466 51940 5485 51996
rect 5541 51940 5560 51996
rect 5466 51912 5560 51940
rect 8356 52236 8450 52264
rect 8356 52180 8375 52236
rect 8431 52180 8450 52236
rect 8356 52156 8450 52180
rect 8356 52100 8375 52156
rect 8431 52100 8450 52156
rect 8356 52076 8450 52100
rect 8356 52020 8375 52076
rect 8431 52020 8450 52076
rect 8356 51996 8450 52020
rect 8356 51940 8375 51996
rect 8431 51940 8450 51996
rect 8356 51912 8450 51940
rect 11246 52236 11340 52264
rect 11246 52180 11265 52236
rect 11321 52180 11340 52236
rect 11246 52156 11340 52180
rect 11246 52100 11265 52156
rect 11321 52100 11340 52156
rect 11246 52076 11340 52100
rect 11246 52020 11265 52076
rect 11321 52020 11340 52076
rect 11246 51996 11340 52020
rect 11246 51940 11265 51996
rect 11321 51940 11340 51996
rect 11246 51912 11340 51940
rect 14136 52236 14230 52264
rect 14136 52180 14155 52236
rect 14211 52180 14230 52236
rect 14136 52156 14230 52180
rect 14136 52100 14155 52156
rect 14211 52100 14230 52156
rect 14136 52076 14230 52100
rect 14136 52020 14155 52076
rect 14211 52020 14230 52076
rect 14136 51996 14230 52020
rect 14136 51940 14155 51996
rect 14211 51940 14230 51996
rect 14136 51912 14230 51940
rect 17026 52236 17120 52264
rect 17026 52180 17045 52236
rect 17101 52180 17120 52236
rect 17026 52156 17120 52180
rect 17026 52100 17045 52156
rect 17101 52100 17120 52156
rect 17026 52076 17120 52100
rect 17026 52020 17045 52076
rect 17101 52020 17120 52076
rect 17026 51996 17120 52020
rect 17026 51940 17045 51996
rect 17101 51940 17120 51996
rect 17026 51912 17120 51940
rect 19916 52236 20010 52264
rect 19916 52180 19935 52236
rect 19991 52180 20010 52236
rect 19916 52156 20010 52180
rect 19916 52100 19935 52156
rect 19991 52100 20010 52156
rect 19916 52076 20010 52100
rect 19916 52020 19935 52076
rect 19991 52020 20010 52076
rect 19916 51996 20010 52020
rect 19916 51940 19935 51996
rect 19991 51940 20010 51996
rect 19916 51912 20010 51940
rect 22806 52236 22900 52264
rect 22806 52180 22825 52236
rect 22881 52180 22900 52236
rect 22806 52156 22900 52180
rect 22806 52100 22825 52156
rect 22881 52100 22900 52156
rect 22806 52076 22900 52100
rect 22806 52020 22825 52076
rect 22881 52020 22900 52076
rect 22806 51996 22900 52020
rect 22806 51940 22825 51996
rect 22881 51940 22900 51996
rect 22806 51912 22900 51940
rect 25696 52236 25790 52264
rect 25696 52180 25715 52236
rect 25771 52180 25790 52236
rect 25696 52156 25790 52180
rect 25696 52100 25715 52156
rect 25771 52100 25790 52156
rect 25696 52076 25790 52100
rect 25696 52020 25715 52076
rect 25771 52020 25790 52076
rect 25696 51996 25790 52020
rect 25696 51940 25715 51996
rect 25771 51940 25790 51996
rect 25696 51912 25790 51940
rect 28586 52236 28680 52264
rect 28586 52180 28605 52236
rect 28661 52180 28680 52236
rect 28586 52156 28680 52180
rect 28586 52100 28605 52156
rect 28661 52100 28680 52156
rect 28586 52076 28680 52100
rect 28586 52020 28605 52076
rect 28661 52020 28680 52076
rect 28586 51996 28680 52020
rect 28586 51940 28605 51996
rect 28661 51940 28680 51996
rect 28586 51912 28680 51940
rect 31476 52236 31570 52264
rect 31476 52180 31495 52236
rect 31551 52180 31570 52236
rect 31476 52156 31570 52180
rect 31476 52100 31495 52156
rect 31551 52100 31570 52156
rect 31476 52076 31570 52100
rect 31476 52020 31495 52076
rect 31551 52020 31570 52076
rect 31476 51996 31570 52020
rect 31476 51940 31495 51996
rect 31551 51940 31570 51996
rect 31476 51912 31570 51940
rect 34366 52236 34460 52264
rect 34366 52180 34385 52236
rect 34441 52180 34460 52236
rect 34366 52156 34460 52180
rect 34366 52100 34385 52156
rect 34441 52100 34460 52156
rect 34366 52076 34460 52100
rect 34366 52020 34385 52076
rect 34441 52020 34460 52076
rect 34366 51996 34460 52020
rect 34366 51940 34385 51996
rect 34441 51940 34460 51996
rect 34366 51912 34460 51940
rect 37256 52236 37350 52264
rect 37256 52180 37275 52236
rect 37331 52180 37350 52236
rect 37256 52156 37350 52180
rect 37256 52100 37275 52156
rect 37331 52100 37350 52156
rect 37256 52076 37350 52100
rect 37256 52020 37275 52076
rect 37331 52020 37350 52076
rect 37256 51996 37350 52020
rect 37256 51940 37275 51996
rect 37331 51940 37350 51996
rect 37256 51912 37350 51940
rect 40146 52236 40240 52264
rect 40146 52180 40165 52236
rect 40221 52180 40240 52236
rect 40146 52156 40240 52180
rect 40146 52100 40165 52156
rect 40221 52100 40240 52156
rect 40146 52076 40240 52100
rect 40146 52020 40165 52076
rect 40221 52020 40240 52076
rect 40146 51996 40240 52020
rect 40146 51940 40165 51996
rect 40221 51940 40240 51996
rect 40146 51912 40240 51940
rect 43036 52236 43130 52264
rect 43036 52180 43055 52236
rect 43111 52180 43130 52236
rect 43036 52156 43130 52180
rect 43036 52100 43055 52156
rect 43111 52100 43130 52156
rect 43036 52076 43130 52100
rect 43036 52020 43055 52076
rect 43111 52020 43130 52076
rect 43036 51996 43130 52020
rect 43036 51940 43055 51996
rect 43111 51940 43130 51996
rect 43036 51912 43130 51940
rect 45926 52236 46020 52264
rect 45926 52180 45945 52236
rect 46001 52180 46020 52236
rect 45926 52156 46020 52180
rect 45926 52100 45945 52156
rect 46001 52100 46020 52156
rect 45926 52076 46020 52100
rect 45926 52020 45945 52076
rect 46001 52020 46020 52076
rect 45926 51996 46020 52020
rect 45926 51940 45945 51996
rect 46001 51940 46020 51996
rect 45926 51912 46020 51940
rect 48873 52236 48967 52264
rect 48873 52180 48892 52236
rect 48948 52180 48967 52236
rect 48873 52156 48967 52180
rect 48873 52100 48892 52156
rect 48948 52100 48967 52156
rect 48873 52076 48967 52100
rect 48873 52020 48892 52076
rect 48948 52020 48967 52076
rect 48873 51996 48967 52020
rect 48873 51940 48892 51996
rect 48948 51940 48967 51996
rect 48873 51912 48967 51940
rect 49722 52236 49922 52264
rect 49722 52180 49754 52236
rect 49810 52180 49834 52236
rect 49890 52180 49922 52236
rect 49722 52156 49922 52180
rect 49722 52100 49754 52156
rect 49810 52100 49834 52156
rect 49890 52100 49922 52156
rect 49722 52076 49922 52100
rect 49722 52020 49754 52076
rect 49810 52020 49834 52076
rect 49890 52020 49922 52076
rect 49722 51996 49922 52020
rect 49722 51940 49754 51996
rect 49810 51940 49834 51996
rect 49890 51940 49922 51996
rect 49722 51912 49922 51940
rect 53012 52236 53140 52264
rect 53012 52180 53048 52236
rect 53104 52180 53140 52236
rect 53012 52156 53140 52180
rect 53012 52100 53048 52156
rect 53104 52100 53140 52156
rect 53012 52076 53140 52100
rect 53012 52020 53048 52076
rect 53104 52020 53140 52076
rect 53012 51996 53140 52020
rect 53012 51940 53048 51996
rect 53104 51940 53140 51996
rect 53012 51912 53140 51940
rect 53170 52236 53298 52264
rect 53170 52180 53206 52236
rect 53262 52180 53298 52236
rect 53170 52156 53298 52180
rect 53170 52100 53206 52156
rect 53262 52100 53298 52156
rect 53170 52076 53298 52100
rect 53170 52020 53206 52076
rect 53262 52020 53298 52076
rect 53170 51996 53298 52020
rect 53170 51940 53206 51996
rect 53262 51940 53298 51996
rect 53170 51912 53298 51940
rect 53526 52236 53654 52264
rect 53526 52180 53562 52236
rect 53618 52180 53654 52236
rect 53526 52156 53654 52180
rect 53526 52100 53562 52156
rect 53618 52100 53654 52156
rect 53526 52076 53654 52100
rect 53526 52020 53562 52076
rect 53618 52020 53654 52076
rect 53526 51996 53654 52020
rect 53526 51940 53562 51996
rect 53618 51940 53654 51996
rect 53526 51912 53654 51940
rect 54844 52236 54972 52264
rect 54844 52180 54880 52236
rect 54936 52180 54972 52236
rect 54844 52156 54972 52180
rect 54844 52100 54880 52156
rect 54936 52100 54972 52156
rect 54844 52076 54972 52100
rect 54844 52020 54880 52076
rect 54936 52020 54972 52076
rect 54844 51996 54972 52020
rect 54844 51940 54880 51996
rect 54936 51940 54972 51996
rect 54844 51912 54972 51940
rect 55437 52236 55565 52264
rect 55437 52180 55473 52236
rect 55529 52180 55565 52236
rect 55437 52156 55565 52180
rect 55437 52100 55473 52156
rect 55529 52100 55565 52156
rect 55437 52076 55565 52100
rect 55437 52020 55473 52076
rect 55529 52020 55565 52076
rect 55437 51996 55565 52020
rect 55437 51940 55473 51996
rect 55529 51940 55565 51996
rect 55437 51912 55565 51940
rect 56583 52236 56711 52264
rect 56583 52180 56619 52236
rect 56675 52180 56711 52236
rect 56583 52156 56711 52180
rect 56583 52100 56619 52156
rect 56675 52100 56711 52156
rect 56583 52076 56711 52100
rect 56583 52020 56619 52076
rect 56675 52020 56711 52076
rect 56583 51996 56711 52020
rect 56583 51940 56619 51996
rect 56675 51940 56711 51996
rect 56583 51912 56711 51940
rect 58033 52236 58213 52264
rect 58033 52180 58055 52236
rect 58111 52180 58135 52236
rect 58191 52180 58213 52236
rect 58033 52156 58213 52180
rect 58033 52100 58055 52156
rect 58111 52100 58135 52156
rect 58191 52100 58213 52156
rect 58033 52076 58213 52100
rect 58033 52020 58055 52076
rect 58111 52020 58135 52076
rect 58191 52020 58213 52076
rect 58033 51996 58213 52020
rect 58033 51940 58055 51996
rect 58111 51940 58135 51996
rect 58191 51940 58213 51996
rect 58033 51912 58213 51940
rect 59256 52236 59396 52264
rect 59256 52180 59298 52236
rect 59354 52180 59396 52236
rect 59256 52156 59396 52180
rect 59256 52100 59298 52156
rect 59354 52100 59396 52156
rect 59256 52076 59396 52100
rect 59256 52020 59298 52076
rect 59354 52020 59396 52076
rect 59256 51996 59396 52020
rect 59256 51940 59298 51996
rect 59354 51940 59396 51996
rect 59256 51912 59396 51940
rect 59426 52236 59542 52264
rect 59426 52180 59456 52236
rect 59512 52180 59542 52236
rect 59426 52156 59542 52180
rect 59426 52100 59456 52156
rect 59512 52100 59542 52156
rect 59426 52076 59542 52100
rect 59426 52020 59456 52076
rect 59512 52020 59542 52076
rect 59426 51996 59542 52020
rect 59426 51940 59456 51996
rect 59512 51940 59542 51996
rect 59426 51912 59542 51940
rect 59734 52236 59850 52264
rect 59734 52180 59764 52236
rect 59820 52180 59850 52236
rect 59734 52156 59850 52180
rect 59734 52100 59764 52156
rect 59820 52100 59850 52156
rect 59734 52076 59850 52100
rect 59734 52020 59764 52076
rect 59820 52020 59850 52076
rect 59734 51996 59850 52020
rect 59734 51940 59764 51996
rect 59820 51940 59850 51996
rect 59734 51912 59850 51940
rect 59880 52236 59996 52264
rect 59880 52180 59910 52236
rect 59966 52180 59996 52236
rect 59880 52156 59996 52180
rect 59880 52100 59910 52156
rect 59966 52100 59996 52156
rect 59880 52076 59996 52100
rect 59880 52020 59910 52076
rect 59966 52020 59996 52076
rect 59880 51996 59996 52020
rect 59880 51940 59910 51996
rect 59966 51940 59996 51996
rect 59880 51912 59996 51940
rect 60026 52236 60202 52264
rect 60026 52180 60046 52236
rect 60102 52180 60126 52236
rect 60182 52180 60202 52236
rect 60026 52156 60202 52180
rect 60026 52100 60046 52156
rect 60102 52100 60126 52156
rect 60182 52100 60202 52156
rect 60026 52076 60202 52100
rect 60026 52020 60046 52076
rect 60102 52020 60126 52076
rect 60182 52020 60202 52076
rect 60026 51996 60202 52020
rect 60026 51940 60046 51996
rect 60102 51940 60126 51996
rect 60182 51940 60202 51996
rect 60026 51912 60202 51940
rect 62399 52236 62573 52264
rect 62399 52180 62418 52236
rect 62474 52180 62498 52236
rect 62554 52180 62573 52236
rect 62399 52156 62573 52180
rect 62399 52100 62418 52156
rect 62474 52100 62498 52156
rect 62554 52100 62573 52156
rect 63512 52126 63540 52566
rect 62399 52076 62573 52100
rect 62399 52020 62418 52076
rect 62474 52020 62498 52076
rect 62554 52020 62573 52076
rect 63500 52120 63552 52126
rect 63500 52062 63552 52068
rect 62399 51996 62573 52020
rect 62399 51940 62418 51996
rect 62474 51940 62498 51996
rect 62554 51940 62573 51996
rect 62399 51912 62573 51940
rect 2112 44588 2216 44616
rect 2112 44532 2136 44588
rect 2192 44532 2216 44588
rect 2112 44508 2216 44532
rect 2112 44452 2136 44508
rect 2192 44452 2216 44508
rect 2112 44428 2216 44452
rect 2112 44372 2136 44428
rect 2192 44372 2216 44428
rect 2112 44348 2216 44372
rect 2112 44292 2136 44348
rect 2192 44292 2216 44348
rect 2112 44264 2216 44292
rect 5613 44588 5707 44616
rect 5613 44532 5632 44588
rect 5688 44532 5707 44588
rect 5613 44508 5707 44532
rect 5613 44452 5632 44508
rect 5688 44452 5707 44508
rect 5613 44428 5707 44452
rect 5613 44372 5632 44428
rect 5688 44372 5707 44428
rect 5613 44348 5707 44372
rect 5613 44292 5632 44348
rect 5688 44292 5707 44348
rect 5613 44264 5707 44292
rect 8503 44588 8597 44616
rect 8503 44532 8522 44588
rect 8578 44532 8597 44588
rect 8503 44508 8597 44532
rect 8503 44452 8522 44508
rect 8578 44452 8597 44508
rect 8503 44428 8597 44452
rect 8503 44372 8522 44428
rect 8578 44372 8597 44428
rect 8503 44348 8597 44372
rect 8503 44292 8522 44348
rect 8578 44292 8597 44348
rect 8503 44264 8597 44292
rect 11393 44588 11487 44616
rect 11393 44532 11412 44588
rect 11468 44532 11487 44588
rect 11393 44508 11487 44532
rect 11393 44452 11412 44508
rect 11468 44452 11487 44508
rect 11393 44428 11487 44452
rect 11393 44372 11412 44428
rect 11468 44372 11487 44428
rect 11393 44348 11487 44372
rect 11393 44292 11412 44348
rect 11468 44292 11487 44348
rect 11393 44264 11487 44292
rect 14283 44588 14377 44616
rect 14283 44532 14302 44588
rect 14358 44532 14377 44588
rect 14283 44508 14377 44532
rect 14283 44452 14302 44508
rect 14358 44452 14377 44508
rect 14283 44428 14377 44452
rect 14283 44372 14302 44428
rect 14358 44372 14377 44428
rect 14283 44348 14377 44372
rect 14283 44292 14302 44348
rect 14358 44292 14377 44348
rect 14283 44264 14377 44292
rect 17173 44588 17267 44616
rect 17173 44532 17192 44588
rect 17248 44532 17267 44588
rect 17173 44508 17267 44532
rect 17173 44452 17192 44508
rect 17248 44452 17267 44508
rect 17173 44428 17267 44452
rect 17173 44372 17192 44428
rect 17248 44372 17267 44428
rect 17173 44348 17267 44372
rect 17173 44292 17192 44348
rect 17248 44292 17267 44348
rect 17173 44264 17267 44292
rect 20063 44588 20157 44616
rect 20063 44532 20082 44588
rect 20138 44532 20157 44588
rect 20063 44508 20157 44532
rect 20063 44452 20082 44508
rect 20138 44452 20157 44508
rect 20063 44428 20157 44452
rect 20063 44372 20082 44428
rect 20138 44372 20157 44428
rect 20063 44348 20157 44372
rect 20063 44292 20082 44348
rect 20138 44292 20157 44348
rect 20063 44264 20157 44292
rect 22953 44588 23047 44616
rect 22953 44532 22972 44588
rect 23028 44532 23047 44588
rect 22953 44508 23047 44532
rect 22953 44452 22972 44508
rect 23028 44452 23047 44508
rect 22953 44428 23047 44452
rect 22953 44372 22972 44428
rect 23028 44372 23047 44428
rect 22953 44348 23047 44372
rect 22953 44292 22972 44348
rect 23028 44292 23047 44348
rect 22953 44264 23047 44292
rect 25843 44588 25937 44616
rect 25843 44532 25862 44588
rect 25918 44532 25937 44588
rect 25843 44508 25937 44532
rect 25843 44452 25862 44508
rect 25918 44452 25937 44508
rect 25843 44428 25937 44452
rect 25843 44372 25862 44428
rect 25918 44372 25937 44428
rect 25843 44348 25937 44372
rect 25843 44292 25862 44348
rect 25918 44292 25937 44348
rect 25843 44264 25937 44292
rect 28733 44588 28827 44616
rect 28733 44532 28752 44588
rect 28808 44532 28827 44588
rect 28733 44508 28827 44532
rect 28733 44452 28752 44508
rect 28808 44452 28827 44508
rect 28733 44428 28827 44452
rect 28733 44372 28752 44428
rect 28808 44372 28827 44428
rect 28733 44348 28827 44372
rect 28733 44292 28752 44348
rect 28808 44292 28827 44348
rect 28733 44264 28827 44292
rect 31623 44588 31717 44616
rect 31623 44532 31642 44588
rect 31698 44532 31717 44588
rect 31623 44508 31717 44532
rect 31623 44452 31642 44508
rect 31698 44452 31717 44508
rect 31623 44428 31717 44452
rect 31623 44372 31642 44428
rect 31698 44372 31717 44428
rect 31623 44348 31717 44372
rect 31623 44292 31642 44348
rect 31698 44292 31717 44348
rect 31623 44264 31717 44292
rect 34513 44588 34607 44616
rect 34513 44532 34532 44588
rect 34588 44532 34607 44588
rect 34513 44508 34607 44532
rect 34513 44452 34532 44508
rect 34588 44452 34607 44508
rect 34513 44428 34607 44452
rect 34513 44372 34532 44428
rect 34588 44372 34607 44428
rect 34513 44348 34607 44372
rect 34513 44292 34532 44348
rect 34588 44292 34607 44348
rect 34513 44264 34607 44292
rect 37403 44588 37497 44616
rect 37403 44532 37422 44588
rect 37478 44532 37497 44588
rect 37403 44508 37497 44532
rect 37403 44452 37422 44508
rect 37478 44452 37497 44508
rect 37403 44428 37497 44452
rect 37403 44372 37422 44428
rect 37478 44372 37497 44428
rect 37403 44348 37497 44372
rect 37403 44292 37422 44348
rect 37478 44292 37497 44348
rect 37403 44264 37497 44292
rect 40293 44588 40387 44616
rect 40293 44532 40312 44588
rect 40368 44532 40387 44588
rect 40293 44508 40387 44532
rect 40293 44452 40312 44508
rect 40368 44452 40387 44508
rect 40293 44428 40387 44452
rect 40293 44372 40312 44428
rect 40368 44372 40387 44428
rect 40293 44348 40387 44372
rect 40293 44292 40312 44348
rect 40368 44292 40387 44348
rect 40293 44264 40387 44292
rect 43183 44588 43277 44616
rect 43183 44532 43202 44588
rect 43258 44532 43277 44588
rect 43183 44508 43277 44532
rect 43183 44452 43202 44508
rect 43258 44452 43277 44508
rect 43183 44428 43277 44452
rect 43183 44372 43202 44428
rect 43258 44372 43277 44428
rect 43183 44348 43277 44372
rect 43183 44292 43202 44348
rect 43258 44292 43277 44348
rect 43183 44264 43277 44292
rect 46073 44588 46167 44616
rect 46073 44532 46092 44588
rect 46148 44532 46167 44588
rect 46073 44508 46167 44532
rect 46073 44452 46092 44508
rect 46148 44452 46167 44508
rect 46073 44428 46167 44452
rect 46073 44372 46092 44428
rect 46148 44372 46167 44428
rect 46073 44348 46167 44372
rect 46073 44292 46092 44348
rect 46148 44292 46167 44348
rect 46073 44264 46167 44292
rect 52302 44588 52412 44616
rect 52302 44532 52329 44588
rect 52385 44532 52412 44588
rect 52302 44508 52412 44532
rect 52302 44452 52329 44508
rect 52385 44452 52412 44508
rect 52302 44428 52412 44452
rect 52302 44372 52329 44428
rect 52385 44372 52412 44428
rect 52302 44348 52412 44372
rect 52302 44292 52329 44348
rect 52385 44292 52412 44348
rect 52302 44264 52412 44292
rect 53694 44588 53822 44616
rect 53694 44532 53730 44588
rect 53786 44532 53822 44588
rect 53694 44508 53822 44532
rect 53694 44452 53730 44508
rect 53786 44452 53822 44508
rect 53694 44428 53822 44452
rect 53694 44372 53730 44428
rect 53786 44372 53822 44428
rect 53694 44348 53822 44372
rect 53694 44292 53730 44348
rect 53786 44292 53822 44348
rect 53694 44264 53822 44292
rect 54606 44588 54734 44616
rect 54606 44532 54642 44588
rect 54698 44532 54734 44588
rect 54606 44508 54734 44532
rect 54606 44452 54642 44508
rect 54698 44452 54734 44508
rect 54606 44428 54734 44452
rect 54606 44372 54642 44428
rect 54698 44372 54734 44428
rect 54606 44348 54734 44372
rect 54606 44292 54642 44348
rect 54698 44292 54734 44348
rect 54606 44264 54734 44292
rect 55002 44588 55118 44616
rect 55002 44532 55032 44588
rect 55088 44532 55118 44588
rect 55002 44508 55118 44532
rect 55002 44452 55032 44508
rect 55088 44452 55118 44508
rect 55002 44428 55118 44452
rect 55002 44372 55032 44428
rect 55088 44372 55118 44428
rect 55002 44348 55118 44372
rect 55002 44292 55032 44348
rect 55088 44292 55118 44348
rect 55002 44264 55118 44292
rect 55712 44588 55840 44616
rect 55712 44532 55748 44588
rect 55804 44532 55840 44588
rect 55712 44508 55840 44532
rect 55712 44452 55748 44508
rect 55804 44452 55840 44508
rect 55712 44428 55840 44452
rect 55712 44372 55748 44428
rect 55804 44372 55840 44428
rect 55712 44348 55840 44372
rect 55712 44292 55748 44348
rect 55804 44292 55840 44348
rect 55712 44264 55840 44292
rect 56290 44588 56418 44616
rect 56290 44532 56326 44588
rect 56382 44532 56418 44588
rect 56290 44508 56418 44532
rect 56290 44452 56326 44508
rect 56382 44452 56418 44508
rect 56290 44428 56418 44452
rect 56290 44372 56326 44428
rect 56382 44372 56418 44428
rect 56290 44348 56418 44372
rect 56290 44292 56326 44348
rect 56382 44292 56418 44348
rect 56290 44264 56418 44292
rect 56741 44588 56857 44616
rect 56741 44532 56771 44588
rect 56827 44532 56857 44588
rect 56741 44508 56857 44532
rect 56741 44452 56771 44508
rect 56827 44452 56857 44508
rect 56741 44428 56857 44452
rect 56741 44372 56771 44428
rect 56827 44372 56857 44428
rect 56741 44348 56857 44372
rect 56741 44292 56771 44348
rect 56827 44292 56857 44348
rect 56741 44264 56857 44292
rect 57045 44588 57161 44616
rect 57045 44532 57075 44588
rect 57131 44532 57161 44588
rect 57045 44508 57161 44532
rect 57045 44452 57075 44508
rect 57131 44452 57161 44508
rect 57045 44428 57161 44452
rect 57045 44372 57075 44428
rect 57131 44372 57161 44428
rect 57045 44348 57161 44372
rect 57045 44292 57075 44348
rect 57131 44292 57161 44348
rect 57045 44264 57161 44292
rect 57887 44588 58003 44616
rect 57887 44532 57917 44588
rect 57973 44532 58003 44588
rect 57887 44508 58003 44532
rect 57887 44452 57917 44508
rect 57973 44452 58003 44508
rect 57887 44428 58003 44452
rect 57887 44372 57917 44428
rect 57973 44372 58003 44428
rect 57887 44348 58003 44372
rect 57887 44292 57917 44348
rect 57973 44292 58003 44348
rect 57887 44264 58003 44292
rect 58437 44588 58501 44616
rect 58437 44532 58441 44588
rect 58497 44532 58501 44588
rect 58437 44508 58501 44532
rect 58437 44452 58441 44508
rect 58497 44452 58501 44508
rect 58437 44428 58501 44452
rect 58437 44372 58441 44428
rect 58497 44372 58501 44428
rect 58437 44348 58501 44372
rect 58437 44292 58441 44348
rect 58497 44292 58501 44348
rect 58437 44264 58501 44292
rect 59110 44588 59226 44616
rect 59110 44532 59140 44588
rect 59196 44532 59226 44588
rect 59110 44508 59226 44532
rect 59110 44452 59140 44508
rect 59196 44452 59226 44508
rect 59110 44428 59226 44452
rect 59110 44372 59140 44428
rect 59196 44372 59226 44428
rect 59110 44348 59226 44372
rect 59110 44292 59140 44348
rect 59196 44292 59226 44348
rect 59110 44264 59226 44292
rect 60388 44588 60504 44616
rect 60388 44532 60418 44588
rect 60474 44532 60504 44588
rect 60388 44508 60504 44532
rect 60388 44452 60418 44508
rect 60474 44452 60504 44508
rect 60388 44428 60504 44452
rect 60388 44372 60418 44428
rect 60474 44372 60504 44428
rect 60388 44348 60504 44372
rect 60388 44292 60418 44348
rect 60474 44292 60504 44348
rect 60388 44264 60504 44292
rect 60546 44588 60662 44616
rect 60546 44532 60576 44588
rect 60632 44532 60662 44588
rect 60546 44508 60662 44532
rect 60546 44452 60576 44508
rect 60632 44452 60662 44508
rect 60546 44428 60662 44452
rect 60546 44372 60576 44428
rect 60632 44372 60662 44428
rect 60546 44348 60662 44372
rect 60546 44292 60576 44348
rect 60632 44292 60662 44348
rect 60546 44264 60662 44292
rect 62601 44588 62775 44616
rect 62601 44532 62620 44588
rect 62676 44532 62700 44588
rect 62756 44532 62775 44588
rect 62601 44508 62775 44532
rect 62601 44452 62620 44508
rect 62676 44452 62700 44508
rect 62756 44452 62775 44508
rect 62601 44428 62775 44452
rect 62601 44372 62620 44428
rect 62676 44372 62700 44428
rect 62756 44372 62775 44428
rect 62601 44348 62775 44372
rect 62601 44292 62620 44348
rect 62676 44292 62700 44348
rect 62756 44292 62775 44348
rect 62601 44264 62775 44292
rect 2244 42236 2444 42264
rect 2244 42180 2276 42236
rect 2332 42180 2356 42236
rect 2412 42180 2444 42236
rect 2244 42156 2444 42180
rect 2244 42100 2276 42156
rect 2332 42100 2356 42156
rect 2412 42100 2444 42156
rect 2244 42076 2444 42100
rect 2244 42020 2276 42076
rect 2332 42020 2356 42076
rect 2412 42020 2444 42076
rect 2244 41996 2444 42020
rect 2244 41940 2276 41996
rect 2332 41940 2356 41996
rect 2412 41940 2444 41996
rect 2244 41912 2444 41940
rect 5466 42236 5560 42264
rect 5466 42180 5485 42236
rect 5541 42180 5560 42236
rect 5466 42156 5560 42180
rect 5466 42100 5485 42156
rect 5541 42100 5560 42156
rect 5466 42076 5560 42100
rect 5466 42020 5485 42076
rect 5541 42020 5560 42076
rect 5466 41996 5560 42020
rect 5466 41940 5485 41996
rect 5541 41940 5560 41996
rect 5466 41912 5560 41940
rect 8356 42236 8450 42264
rect 8356 42180 8375 42236
rect 8431 42180 8450 42236
rect 8356 42156 8450 42180
rect 8356 42100 8375 42156
rect 8431 42100 8450 42156
rect 8356 42076 8450 42100
rect 8356 42020 8375 42076
rect 8431 42020 8450 42076
rect 8356 41996 8450 42020
rect 8356 41940 8375 41996
rect 8431 41940 8450 41996
rect 8356 41912 8450 41940
rect 11246 42236 11340 42264
rect 11246 42180 11265 42236
rect 11321 42180 11340 42236
rect 11246 42156 11340 42180
rect 11246 42100 11265 42156
rect 11321 42100 11340 42156
rect 11246 42076 11340 42100
rect 11246 42020 11265 42076
rect 11321 42020 11340 42076
rect 11246 41996 11340 42020
rect 11246 41940 11265 41996
rect 11321 41940 11340 41996
rect 11246 41912 11340 41940
rect 14136 42236 14230 42264
rect 14136 42180 14155 42236
rect 14211 42180 14230 42236
rect 14136 42156 14230 42180
rect 14136 42100 14155 42156
rect 14211 42100 14230 42156
rect 14136 42076 14230 42100
rect 14136 42020 14155 42076
rect 14211 42020 14230 42076
rect 14136 41996 14230 42020
rect 14136 41940 14155 41996
rect 14211 41940 14230 41996
rect 14136 41912 14230 41940
rect 17026 42236 17120 42264
rect 17026 42180 17045 42236
rect 17101 42180 17120 42236
rect 17026 42156 17120 42180
rect 17026 42100 17045 42156
rect 17101 42100 17120 42156
rect 17026 42076 17120 42100
rect 17026 42020 17045 42076
rect 17101 42020 17120 42076
rect 17026 41996 17120 42020
rect 17026 41940 17045 41996
rect 17101 41940 17120 41996
rect 17026 41912 17120 41940
rect 19916 42236 20010 42264
rect 19916 42180 19935 42236
rect 19991 42180 20010 42236
rect 19916 42156 20010 42180
rect 19916 42100 19935 42156
rect 19991 42100 20010 42156
rect 19916 42076 20010 42100
rect 19916 42020 19935 42076
rect 19991 42020 20010 42076
rect 19916 41996 20010 42020
rect 19916 41940 19935 41996
rect 19991 41940 20010 41996
rect 19916 41912 20010 41940
rect 22806 42236 22900 42264
rect 22806 42180 22825 42236
rect 22881 42180 22900 42236
rect 22806 42156 22900 42180
rect 22806 42100 22825 42156
rect 22881 42100 22900 42156
rect 22806 42076 22900 42100
rect 22806 42020 22825 42076
rect 22881 42020 22900 42076
rect 22806 41996 22900 42020
rect 22806 41940 22825 41996
rect 22881 41940 22900 41996
rect 22806 41912 22900 41940
rect 25696 42236 25790 42264
rect 25696 42180 25715 42236
rect 25771 42180 25790 42236
rect 25696 42156 25790 42180
rect 25696 42100 25715 42156
rect 25771 42100 25790 42156
rect 25696 42076 25790 42100
rect 25696 42020 25715 42076
rect 25771 42020 25790 42076
rect 25696 41996 25790 42020
rect 25696 41940 25715 41996
rect 25771 41940 25790 41996
rect 25696 41912 25790 41940
rect 28586 42236 28680 42264
rect 28586 42180 28605 42236
rect 28661 42180 28680 42236
rect 28586 42156 28680 42180
rect 28586 42100 28605 42156
rect 28661 42100 28680 42156
rect 28586 42076 28680 42100
rect 28586 42020 28605 42076
rect 28661 42020 28680 42076
rect 28586 41996 28680 42020
rect 28586 41940 28605 41996
rect 28661 41940 28680 41996
rect 28586 41912 28680 41940
rect 31476 42236 31570 42264
rect 31476 42180 31495 42236
rect 31551 42180 31570 42236
rect 31476 42156 31570 42180
rect 31476 42100 31495 42156
rect 31551 42100 31570 42156
rect 31476 42076 31570 42100
rect 31476 42020 31495 42076
rect 31551 42020 31570 42076
rect 31476 41996 31570 42020
rect 31476 41940 31495 41996
rect 31551 41940 31570 41996
rect 31476 41912 31570 41940
rect 34366 42236 34460 42264
rect 34366 42180 34385 42236
rect 34441 42180 34460 42236
rect 34366 42156 34460 42180
rect 34366 42100 34385 42156
rect 34441 42100 34460 42156
rect 34366 42076 34460 42100
rect 34366 42020 34385 42076
rect 34441 42020 34460 42076
rect 34366 41996 34460 42020
rect 34366 41940 34385 41996
rect 34441 41940 34460 41996
rect 34366 41912 34460 41940
rect 37256 42236 37350 42264
rect 37256 42180 37275 42236
rect 37331 42180 37350 42236
rect 37256 42156 37350 42180
rect 37256 42100 37275 42156
rect 37331 42100 37350 42156
rect 37256 42076 37350 42100
rect 37256 42020 37275 42076
rect 37331 42020 37350 42076
rect 37256 41996 37350 42020
rect 37256 41940 37275 41996
rect 37331 41940 37350 41996
rect 37256 41912 37350 41940
rect 40146 42236 40240 42264
rect 40146 42180 40165 42236
rect 40221 42180 40240 42236
rect 40146 42156 40240 42180
rect 40146 42100 40165 42156
rect 40221 42100 40240 42156
rect 40146 42076 40240 42100
rect 40146 42020 40165 42076
rect 40221 42020 40240 42076
rect 40146 41996 40240 42020
rect 40146 41940 40165 41996
rect 40221 41940 40240 41996
rect 40146 41912 40240 41940
rect 43036 42236 43130 42264
rect 43036 42180 43055 42236
rect 43111 42180 43130 42236
rect 43036 42156 43130 42180
rect 43036 42100 43055 42156
rect 43111 42100 43130 42156
rect 43036 42076 43130 42100
rect 43036 42020 43055 42076
rect 43111 42020 43130 42076
rect 43036 41996 43130 42020
rect 43036 41940 43055 41996
rect 43111 41940 43130 41996
rect 43036 41912 43130 41940
rect 45926 42236 46020 42264
rect 45926 42180 45945 42236
rect 46001 42180 46020 42236
rect 45926 42156 46020 42180
rect 45926 42100 45945 42156
rect 46001 42100 46020 42156
rect 45926 42076 46020 42100
rect 45926 42020 45945 42076
rect 46001 42020 46020 42076
rect 45926 41996 46020 42020
rect 45926 41940 45945 41996
rect 46001 41940 46020 41996
rect 45926 41912 46020 41940
rect 48873 42236 48967 42264
rect 48873 42180 48892 42236
rect 48948 42180 48967 42236
rect 48873 42156 48967 42180
rect 48873 42100 48892 42156
rect 48948 42100 48967 42156
rect 48873 42076 48967 42100
rect 48873 42020 48892 42076
rect 48948 42020 48967 42076
rect 48873 41996 48967 42020
rect 48873 41940 48892 41996
rect 48948 41940 48967 41996
rect 48873 41912 48967 41940
rect 49722 42236 49922 42264
rect 49722 42180 49754 42236
rect 49810 42180 49834 42236
rect 49890 42180 49922 42236
rect 49722 42156 49922 42180
rect 49722 42100 49754 42156
rect 49810 42100 49834 42156
rect 49890 42100 49922 42156
rect 49722 42076 49922 42100
rect 49722 42020 49754 42076
rect 49810 42020 49834 42076
rect 49890 42020 49922 42076
rect 49722 41996 49922 42020
rect 49722 41940 49754 41996
rect 49810 41940 49834 41996
rect 49890 41940 49922 41996
rect 49722 41912 49922 41940
rect 53012 42236 53140 42264
rect 53012 42180 53048 42236
rect 53104 42180 53140 42236
rect 53012 42156 53140 42180
rect 53012 42100 53048 42156
rect 53104 42100 53140 42156
rect 53012 42076 53140 42100
rect 53012 42020 53048 42076
rect 53104 42020 53140 42076
rect 53012 41996 53140 42020
rect 53012 41940 53048 41996
rect 53104 41940 53140 41996
rect 53012 41912 53140 41940
rect 53170 42236 53298 42264
rect 53170 42180 53206 42236
rect 53262 42180 53298 42236
rect 53170 42156 53298 42180
rect 53170 42100 53206 42156
rect 53262 42100 53298 42156
rect 53170 42076 53298 42100
rect 53170 42020 53206 42076
rect 53262 42020 53298 42076
rect 53170 41996 53298 42020
rect 53170 41940 53206 41996
rect 53262 41940 53298 41996
rect 53170 41912 53298 41940
rect 53526 42236 53654 42264
rect 53526 42180 53562 42236
rect 53618 42180 53654 42236
rect 53526 42156 53654 42180
rect 53526 42100 53562 42156
rect 53618 42100 53654 42156
rect 53526 42076 53654 42100
rect 53526 42020 53562 42076
rect 53618 42020 53654 42076
rect 53526 41996 53654 42020
rect 53526 41940 53562 41996
rect 53618 41940 53654 41996
rect 53526 41912 53654 41940
rect 54844 42236 54972 42264
rect 54844 42180 54880 42236
rect 54936 42180 54972 42236
rect 54844 42156 54972 42180
rect 54844 42100 54880 42156
rect 54936 42100 54972 42156
rect 54844 42076 54972 42100
rect 54844 42020 54880 42076
rect 54936 42020 54972 42076
rect 54844 41996 54972 42020
rect 54844 41940 54880 41996
rect 54936 41940 54972 41996
rect 54844 41912 54972 41940
rect 55437 42236 55565 42264
rect 55437 42180 55473 42236
rect 55529 42180 55565 42236
rect 55437 42156 55565 42180
rect 55437 42100 55473 42156
rect 55529 42100 55565 42156
rect 55437 42076 55565 42100
rect 55437 42020 55473 42076
rect 55529 42020 55565 42076
rect 55437 41996 55565 42020
rect 55437 41940 55473 41996
rect 55529 41940 55565 41996
rect 55437 41912 55565 41940
rect 56583 42236 56711 42264
rect 56583 42180 56619 42236
rect 56675 42180 56711 42236
rect 56583 42156 56711 42180
rect 56583 42100 56619 42156
rect 56675 42100 56711 42156
rect 56583 42076 56711 42100
rect 56583 42020 56619 42076
rect 56675 42020 56711 42076
rect 56583 41996 56711 42020
rect 56583 41940 56619 41996
rect 56675 41940 56711 41996
rect 56583 41912 56711 41940
rect 58033 42236 58213 42264
rect 58033 42180 58055 42236
rect 58111 42180 58135 42236
rect 58191 42180 58213 42236
rect 58033 42156 58213 42180
rect 58033 42100 58055 42156
rect 58111 42100 58135 42156
rect 58191 42100 58213 42156
rect 58033 42076 58213 42100
rect 58033 42020 58055 42076
rect 58111 42020 58135 42076
rect 58191 42020 58213 42076
rect 58033 41996 58213 42020
rect 58033 41940 58055 41996
rect 58111 41940 58135 41996
rect 58191 41940 58213 41996
rect 58033 41912 58213 41940
rect 59256 42236 59396 42264
rect 59256 42180 59298 42236
rect 59354 42180 59396 42236
rect 59256 42156 59396 42180
rect 59256 42100 59298 42156
rect 59354 42100 59396 42156
rect 59256 42076 59396 42100
rect 59256 42020 59298 42076
rect 59354 42020 59396 42076
rect 59256 41996 59396 42020
rect 59256 41940 59298 41996
rect 59354 41940 59396 41996
rect 59256 41912 59396 41940
rect 59426 42236 59542 42264
rect 59426 42180 59456 42236
rect 59512 42180 59542 42236
rect 59426 42156 59542 42180
rect 59426 42100 59456 42156
rect 59512 42100 59542 42156
rect 59426 42076 59542 42100
rect 59426 42020 59456 42076
rect 59512 42020 59542 42076
rect 59426 41996 59542 42020
rect 59426 41940 59456 41996
rect 59512 41940 59542 41996
rect 59426 41912 59542 41940
rect 59734 42236 59850 42264
rect 59734 42180 59764 42236
rect 59820 42180 59850 42236
rect 59734 42156 59850 42180
rect 59734 42100 59764 42156
rect 59820 42100 59850 42156
rect 59734 42076 59850 42100
rect 59734 42020 59764 42076
rect 59820 42020 59850 42076
rect 59734 41996 59850 42020
rect 59734 41940 59764 41996
rect 59820 41940 59850 41996
rect 59734 41912 59850 41940
rect 59880 42236 59996 42264
rect 59880 42180 59910 42236
rect 59966 42180 59996 42236
rect 59880 42156 59996 42180
rect 59880 42100 59910 42156
rect 59966 42100 59996 42156
rect 59880 42076 59996 42100
rect 59880 42020 59910 42076
rect 59966 42020 59996 42076
rect 59880 41996 59996 42020
rect 59880 41940 59910 41996
rect 59966 41940 59996 41996
rect 59880 41912 59996 41940
rect 60026 42236 60202 42264
rect 60026 42180 60046 42236
rect 60102 42180 60126 42236
rect 60182 42180 60202 42236
rect 60026 42156 60202 42180
rect 60026 42100 60046 42156
rect 60102 42100 60126 42156
rect 60182 42100 60202 42156
rect 60026 42076 60202 42100
rect 60026 42020 60046 42076
rect 60102 42020 60126 42076
rect 60182 42020 60202 42076
rect 60026 41996 60202 42020
rect 60026 41940 60046 41996
rect 60102 41940 60126 41996
rect 60182 41940 60202 41996
rect 60026 41912 60202 41940
rect 62399 42236 62573 42264
rect 62399 42180 62418 42236
rect 62474 42180 62498 42236
rect 62554 42180 62573 42236
rect 62399 42156 62573 42180
rect 62399 42100 62418 42156
rect 62474 42100 62498 42156
rect 62554 42100 62573 42156
rect 62399 42076 62573 42100
rect 62399 42020 62418 42076
rect 62474 42020 62498 42076
rect 62554 42020 62573 42076
rect 62399 41996 62573 42020
rect 62399 41940 62418 41996
rect 62474 41940 62498 41996
rect 62554 41940 62573 41996
rect 62399 41912 62573 41940
rect 63500 41744 63552 41750
rect 63500 41686 63552 41692
rect 63512 39574 63540 41686
rect 63500 39568 63552 39574
rect 63500 39510 63552 39516
rect 63512 38010 63540 39510
rect 63500 38004 63552 38010
rect 63500 37946 63552 37952
rect 63500 37868 63552 37874
rect 63500 37810 63552 37816
rect 2112 34588 2216 34616
rect 2112 34532 2136 34588
rect 2192 34532 2216 34588
rect 2112 34508 2216 34532
rect 2112 34452 2136 34508
rect 2192 34452 2216 34508
rect 2112 34428 2216 34452
rect 2112 34372 2136 34428
rect 2192 34372 2216 34428
rect 2112 34348 2216 34372
rect 2112 34292 2136 34348
rect 2192 34292 2216 34348
rect 2112 34264 2216 34292
rect 5613 34588 5707 34616
rect 5613 34532 5632 34588
rect 5688 34532 5707 34588
rect 5613 34508 5707 34532
rect 5613 34452 5632 34508
rect 5688 34452 5707 34508
rect 5613 34428 5707 34452
rect 5613 34372 5632 34428
rect 5688 34372 5707 34428
rect 5613 34348 5707 34372
rect 5613 34292 5632 34348
rect 5688 34292 5707 34348
rect 5613 34264 5707 34292
rect 8503 34588 8597 34616
rect 8503 34532 8522 34588
rect 8578 34532 8597 34588
rect 8503 34508 8597 34532
rect 8503 34452 8522 34508
rect 8578 34452 8597 34508
rect 8503 34428 8597 34452
rect 8503 34372 8522 34428
rect 8578 34372 8597 34428
rect 8503 34348 8597 34372
rect 8503 34292 8522 34348
rect 8578 34292 8597 34348
rect 8503 34264 8597 34292
rect 11393 34588 11487 34616
rect 11393 34532 11412 34588
rect 11468 34532 11487 34588
rect 11393 34508 11487 34532
rect 11393 34452 11412 34508
rect 11468 34452 11487 34508
rect 11393 34428 11487 34452
rect 11393 34372 11412 34428
rect 11468 34372 11487 34428
rect 11393 34348 11487 34372
rect 11393 34292 11412 34348
rect 11468 34292 11487 34348
rect 11393 34264 11487 34292
rect 14283 34588 14377 34616
rect 14283 34532 14302 34588
rect 14358 34532 14377 34588
rect 14283 34508 14377 34532
rect 14283 34452 14302 34508
rect 14358 34452 14377 34508
rect 14283 34428 14377 34452
rect 14283 34372 14302 34428
rect 14358 34372 14377 34428
rect 14283 34348 14377 34372
rect 14283 34292 14302 34348
rect 14358 34292 14377 34348
rect 14283 34264 14377 34292
rect 17173 34588 17267 34616
rect 17173 34532 17192 34588
rect 17248 34532 17267 34588
rect 17173 34508 17267 34532
rect 17173 34452 17192 34508
rect 17248 34452 17267 34508
rect 17173 34428 17267 34452
rect 17173 34372 17192 34428
rect 17248 34372 17267 34428
rect 17173 34348 17267 34372
rect 17173 34292 17192 34348
rect 17248 34292 17267 34348
rect 17173 34264 17267 34292
rect 20063 34588 20157 34616
rect 20063 34532 20082 34588
rect 20138 34532 20157 34588
rect 20063 34508 20157 34532
rect 20063 34452 20082 34508
rect 20138 34452 20157 34508
rect 20063 34428 20157 34452
rect 20063 34372 20082 34428
rect 20138 34372 20157 34428
rect 20063 34348 20157 34372
rect 20063 34292 20082 34348
rect 20138 34292 20157 34348
rect 20063 34264 20157 34292
rect 22953 34588 23047 34616
rect 22953 34532 22972 34588
rect 23028 34532 23047 34588
rect 22953 34508 23047 34532
rect 22953 34452 22972 34508
rect 23028 34452 23047 34508
rect 22953 34428 23047 34452
rect 22953 34372 22972 34428
rect 23028 34372 23047 34428
rect 22953 34348 23047 34372
rect 22953 34292 22972 34348
rect 23028 34292 23047 34348
rect 22953 34264 23047 34292
rect 25843 34588 25937 34616
rect 25843 34532 25862 34588
rect 25918 34532 25937 34588
rect 25843 34508 25937 34532
rect 25843 34452 25862 34508
rect 25918 34452 25937 34508
rect 25843 34428 25937 34452
rect 25843 34372 25862 34428
rect 25918 34372 25937 34428
rect 25843 34348 25937 34372
rect 25843 34292 25862 34348
rect 25918 34292 25937 34348
rect 25843 34264 25937 34292
rect 28733 34588 28827 34616
rect 28733 34532 28752 34588
rect 28808 34532 28827 34588
rect 28733 34508 28827 34532
rect 28733 34452 28752 34508
rect 28808 34452 28827 34508
rect 28733 34428 28827 34452
rect 28733 34372 28752 34428
rect 28808 34372 28827 34428
rect 28733 34348 28827 34372
rect 28733 34292 28752 34348
rect 28808 34292 28827 34348
rect 28733 34264 28827 34292
rect 31623 34588 31717 34616
rect 31623 34532 31642 34588
rect 31698 34532 31717 34588
rect 31623 34508 31717 34532
rect 31623 34452 31642 34508
rect 31698 34452 31717 34508
rect 31623 34428 31717 34452
rect 31623 34372 31642 34428
rect 31698 34372 31717 34428
rect 31623 34348 31717 34372
rect 31623 34292 31642 34348
rect 31698 34292 31717 34348
rect 31623 34264 31717 34292
rect 34513 34588 34607 34616
rect 34513 34532 34532 34588
rect 34588 34532 34607 34588
rect 34513 34508 34607 34532
rect 34513 34452 34532 34508
rect 34588 34452 34607 34508
rect 34513 34428 34607 34452
rect 34513 34372 34532 34428
rect 34588 34372 34607 34428
rect 34513 34348 34607 34372
rect 34513 34292 34532 34348
rect 34588 34292 34607 34348
rect 34513 34264 34607 34292
rect 37403 34588 37497 34616
rect 37403 34532 37422 34588
rect 37478 34532 37497 34588
rect 37403 34508 37497 34532
rect 37403 34452 37422 34508
rect 37478 34452 37497 34508
rect 37403 34428 37497 34452
rect 37403 34372 37422 34428
rect 37478 34372 37497 34428
rect 37403 34348 37497 34372
rect 37403 34292 37422 34348
rect 37478 34292 37497 34348
rect 37403 34264 37497 34292
rect 40293 34588 40387 34616
rect 40293 34532 40312 34588
rect 40368 34532 40387 34588
rect 40293 34508 40387 34532
rect 40293 34452 40312 34508
rect 40368 34452 40387 34508
rect 40293 34428 40387 34452
rect 40293 34372 40312 34428
rect 40368 34372 40387 34428
rect 40293 34348 40387 34372
rect 40293 34292 40312 34348
rect 40368 34292 40387 34348
rect 40293 34264 40387 34292
rect 43183 34588 43277 34616
rect 43183 34532 43202 34588
rect 43258 34532 43277 34588
rect 43183 34508 43277 34532
rect 43183 34452 43202 34508
rect 43258 34452 43277 34508
rect 43183 34428 43277 34452
rect 43183 34372 43202 34428
rect 43258 34372 43277 34428
rect 43183 34348 43277 34372
rect 43183 34292 43202 34348
rect 43258 34292 43277 34348
rect 43183 34264 43277 34292
rect 46073 34588 46167 34616
rect 46073 34532 46092 34588
rect 46148 34532 46167 34588
rect 46073 34508 46167 34532
rect 46073 34452 46092 34508
rect 46148 34452 46167 34508
rect 46073 34428 46167 34452
rect 46073 34372 46092 34428
rect 46148 34372 46167 34428
rect 46073 34348 46167 34372
rect 46073 34292 46092 34348
rect 46148 34292 46167 34348
rect 46073 34264 46167 34292
rect 49081 34588 49175 34616
rect 49081 34532 49100 34588
rect 49156 34532 49175 34588
rect 49081 34508 49175 34532
rect 49081 34452 49100 34508
rect 49156 34452 49175 34508
rect 49081 34428 49175 34452
rect 49081 34372 49100 34428
rect 49156 34372 49175 34428
rect 49081 34348 49175 34372
rect 49081 34292 49100 34348
rect 49156 34292 49175 34348
rect 49081 34264 49175 34292
rect 52302 34588 52412 34616
rect 52302 34532 52329 34588
rect 52385 34532 52412 34588
rect 52302 34508 52412 34532
rect 52302 34452 52329 34508
rect 52385 34452 52412 34508
rect 52302 34428 52412 34452
rect 52302 34372 52329 34428
rect 52385 34372 52412 34428
rect 52302 34348 52412 34372
rect 52302 34292 52329 34348
rect 52385 34292 52412 34348
rect 52302 34264 52412 34292
rect 53694 34588 53822 34616
rect 53694 34532 53730 34588
rect 53786 34532 53822 34588
rect 53694 34508 53822 34532
rect 53694 34452 53730 34508
rect 53786 34452 53822 34508
rect 53694 34428 53822 34452
rect 53694 34372 53730 34428
rect 53786 34372 53822 34428
rect 53694 34348 53822 34372
rect 53694 34292 53730 34348
rect 53786 34292 53822 34348
rect 53694 34264 53822 34292
rect 53862 34588 53990 34616
rect 53862 34532 53898 34588
rect 53954 34532 53990 34588
rect 53862 34508 53990 34532
rect 53862 34452 53898 34508
rect 53954 34452 53990 34508
rect 53862 34428 53990 34452
rect 53862 34372 53898 34428
rect 53954 34372 53990 34428
rect 53862 34348 53990 34372
rect 53862 34292 53898 34348
rect 53954 34292 53990 34348
rect 53862 34264 53990 34292
rect 54606 34588 54734 34616
rect 54606 34532 54642 34588
rect 54698 34532 54734 34588
rect 54606 34508 54734 34532
rect 54606 34452 54642 34508
rect 54698 34452 54734 34508
rect 54606 34428 54734 34452
rect 54606 34372 54642 34428
rect 54698 34372 54734 34428
rect 54606 34348 54734 34372
rect 54606 34292 54642 34348
rect 54698 34292 54734 34348
rect 54606 34264 54734 34292
rect 55002 34588 55118 34616
rect 55002 34532 55032 34588
rect 55088 34532 55118 34588
rect 55002 34508 55118 34532
rect 55002 34452 55032 34508
rect 55088 34452 55118 34508
rect 55002 34428 55118 34452
rect 55002 34372 55032 34428
rect 55088 34372 55118 34428
rect 55002 34348 55118 34372
rect 55002 34292 55032 34348
rect 55088 34292 55118 34348
rect 55002 34264 55118 34292
rect 55712 34588 55840 34616
rect 55712 34532 55748 34588
rect 55804 34532 55840 34588
rect 55712 34508 55840 34532
rect 55712 34452 55748 34508
rect 55804 34452 55840 34508
rect 55712 34428 55840 34452
rect 55712 34372 55748 34428
rect 55804 34372 55840 34428
rect 55712 34348 55840 34372
rect 55712 34292 55748 34348
rect 55804 34292 55840 34348
rect 55712 34264 55840 34292
rect 56290 34588 56418 34616
rect 56290 34532 56326 34588
rect 56382 34532 56418 34588
rect 56290 34508 56418 34532
rect 56290 34452 56326 34508
rect 56382 34452 56418 34508
rect 56290 34428 56418 34452
rect 56290 34372 56326 34428
rect 56382 34372 56418 34428
rect 56290 34348 56418 34372
rect 56290 34292 56326 34348
rect 56382 34292 56418 34348
rect 56290 34264 56418 34292
rect 56741 34588 56857 34616
rect 56741 34532 56771 34588
rect 56827 34532 56857 34588
rect 56741 34508 56857 34532
rect 56741 34452 56771 34508
rect 56827 34452 56857 34508
rect 56741 34428 56857 34452
rect 56741 34372 56771 34428
rect 56827 34372 56857 34428
rect 56741 34348 56857 34372
rect 56741 34292 56771 34348
rect 56827 34292 56857 34348
rect 56741 34264 56857 34292
rect 57045 34588 57161 34616
rect 57045 34532 57075 34588
rect 57131 34532 57161 34588
rect 57045 34508 57161 34532
rect 57045 34452 57075 34508
rect 57131 34452 57161 34508
rect 57045 34428 57161 34452
rect 57045 34372 57075 34428
rect 57131 34372 57161 34428
rect 57045 34348 57161 34372
rect 57045 34292 57075 34348
rect 57131 34292 57161 34348
rect 57045 34264 57161 34292
rect 57887 34588 58003 34616
rect 57887 34532 57917 34588
rect 57973 34532 58003 34588
rect 57887 34508 58003 34532
rect 57887 34452 57917 34508
rect 57973 34452 58003 34508
rect 57887 34428 58003 34452
rect 57887 34372 57917 34428
rect 57973 34372 58003 34428
rect 57887 34348 58003 34372
rect 57887 34292 57917 34348
rect 57973 34292 58003 34348
rect 57887 34264 58003 34292
rect 58553 34588 58617 34616
rect 58553 34532 58557 34588
rect 58613 34532 58617 34588
rect 58553 34508 58617 34532
rect 58553 34452 58557 34508
rect 58613 34452 58617 34508
rect 58553 34428 58617 34452
rect 58553 34372 58557 34428
rect 58613 34372 58617 34428
rect 58553 34348 58617 34372
rect 58553 34292 58557 34348
rect 58613 34292 58617 34348
rect 58553 34264 58617 34292
rect 59110 34588 59226 34616
rect 59110 34532 59140 34588
rect 59196 34532 59226 34588
rect 59110 34508 59226 34532
rect 59110 34452 59140 34508
rect 59196 34452 59226 34508
rect 59110 34428 59226 34452
rect 59110 34372 59140 34428
rect 59196 34372 59226 34428
rect 59110 34348 59226 34372
rect 59110 34292 59140 34348
rect 59196 34292 59226 34348
rect 59110 34264 59226 34292
rect 60388 34588 60504 34616
rect 60388 34532 60418 34588
rect 60474 34532 60504 34588
rect 60388 34508 60504 34532
rect 60388 34452 60418 34508
rect 60474 34452 60504 34508
rect 60388 34428 60504 34452
rect 60388 34372 60418 34428
rect 60474 34372 60504 34428
rect 60388 34348 60504 34372
rect 60388 34292 60418 34348
rect 60474 34292 60504 34348
rect 60388 34264 60504 34292
rect 60546 34588 60662 34616
rect 60546 34532 60576 34588
rect 60632 34532 60662 34588
rect 60546 34508 60662 34532
rect 60546 34452 60576 34508
rect 60632 34452 60662 34508
rect 60546 34428 60662 34452
rect 60546 34372 60576 34428
rect 60632 34372 60662 34428
rect 60546 34348 60662 34372
rect 60546 34292 60576 34348
rect 60632 34292 60662 34348
rect 60546 34264 60662 34292
rect 62601 34588 62775 34616
rect 62601 34532 62620 34588
rect 62676 34532 62700 34588
rect 62756 34532 62775 34588
rect 62601 34508 62775 34532
rect 62601 34452 62620 34508
rect 62676 34452 62700 34508
rect 62756 34452 62775 34508
rect 62601 34428 62775 34452
rect 62601 34372 62620 34428
rect 62676 34372 62700 34428
rect 62756 34372 62775 34428
rect 62601 34348 62775 34372
rect 62601 34292 62620 34348
rect 62676 34292 62700 34348
rect 62756 34292 62775 34348
rect 62601 34264 62775 34292
rect 2244 32236 2444 32264
rect 2244 32180 2276 32236
rect 2332 32180 2356 32236
rect 2412 32180 2444 32236
rect 2244 32156 2444 32180
rect 2244 32100 2276 32156
rect 2332 32100 2356 32156
rect 2412 32100 2444 32156
rect 2244 32076 2444 32100
rect 2244 32020 2276 32076
rect 2332 32020 2356 32076
rect 2412 32020 2444 32076
rect 2244 31996 2444 32020
rect 2244 31940 2276 31996
rect 2332 31940 2356 31996
rect 2412 31940 2444 31996
rect 2244 31912 2444 31940
rect 5466 32236 5560 32264
rect 5466 32180 5485 32236
rect 5541 32180 5560 32236
rect 5466 32156 5560 32180
rect 5466 32100 5485 32156
rect 5541 32100 5560 32156
rect 5466 32076 5560 32100
rect 5466 32020 5485 32076
rect 5541 32020 5560 32076
rect 5466 31996 5560 32020
rect 5466 31940 5485 31996
rect 5541 31940 5560 31996
rect 5466 31912 5560 31940
rect 8356 32236 8450 32264
rect 8356 32180 8375 32236
rect 8431 32180 8450 32236
rect 8356 32156 8450 32180
rect 8356 32100 8375 32156
rect 8431 32100 8450 32156
rect 8356 32076 8450 32100
rect 8356 32020 8375 32076
rect 8431 32020 8450 32076
rect 8356 31996 8450 32020
rect 8356 31940 8375 31996
rect 8431 31940 8450 31996
rect 8356 31912 8450 31940
rect 11246 32236 11340 32264
rect 11246 32180 11265 32236
rect 11321 32180 11340 32236
rect 11246 32156 11340 32180
rect 11246 32100 11265 32156
rect 11321 32100 11340 32156
rect 11246 32076 11340 32100
rect 11246 32020 11265 32076
rect 11321 32020 11340 32076
rect 11246 31996 11340 32020
rect 11246 31940 11265 31996
rect 11321 31940 11340 31996
rect 11246 31912 11340 31940
rect 14136 32236 14230 32264
rect 14136 32180 14155 32236
rect 14211 32180 14230 32236
rect 14136 32156 14230 32180
rect 14136 32100 14155 32156
rect 14211 32100 14230 32156
rect 14136 32076 14230 32100
rect 14136 32020 14155 32076
rect 14211 32020 14230 32076
rect 14136 31996 14230 32020
rect 14136 31940 14155 31996
rect 14211 31940 14230 31996
rect 14136 31912 14230 31940
rect 17026 32236 17120 32264
rect 17026 32180 17045 32236
rect 17101 32180 17120 32236
rect 17026 32156 17120 32180
rect 17026 32100 17045 32156
rect 17101 32100 17120 32156
rect 17026 32076 17120 32100
rect 17026 32020 17045 32076
rect 17101 32020 17120 32076
rect 17026 31996 17120 32020
rect 17026 31940 17045 31996
rect 17101 31940 17120 31996
rect 17026 31912 17120 31940
rect 19916 32236 20010 32264
rect 19916 32180 19935 32236
rect 19991 32180 20010 32236
rect 19916 32156 20010 32180
rect 19916 32100 19935 32156
rect 19991 32100 20010 32156
rect 19916 32076 20010 32100
rect 19916 32020 19935 32076
rect 19991 32020 20010 32076
rect 19916 31996 20010 32020
rect 19916 31940 19935 31996
rect 19991 31940 20010 31996
rect 19916 31912 20010 31940
rect 22806 32236 22900 32264
rect 22806 32180 22825 32236
rect 22881 32180 22900 32236
rect 22806 32156 22900 32180
rect 22806 32100 22825 32156
rect 22881 32100 22900 32156
rect 22806 32076 22900 32100
rect 22806 32020 22825 32076
rect 22881 32020 22900 32076
rect 22806 31996 22900 32020
rect 22806 31940 22825 31996
rect 22881 31940 22900 31996
rect 22806 31912 22900 31940
rect 25696 32236 25790 32264
rect 25696 32180 25715 32236
rect 25771 32180 25790 32236
rect 25696 32156 25790 32180
rect 25696 32100 25715 32156
rect 25771 32100 25790 32156
rect 25696 32076 25790 32100
rect 25696 32020 25715 32076
rect 25771 32020 25790 32076
rect 25696 31996 25790 32020
rect 25696 31940 25715 31996
rect 25771 31940 25790 31996
rect 25696 31912 25790 31940
rect 28586 32236 28680 32264
rect 28586 32180 28605 32236
rect 28661 32180 28680 32236
rect 28586 32156 28680 32180
rect 28586 32100 28605 32156
rect 28661 32100 28680 32156
rect 28586 32076 28680 32100
rect 28586 32020 28605 32076
rect 28661 32020 28680 32076
rect 28586 31996 28680 32020
rect 28586 31940 28605 31996
rect 28661 31940 28680 31996
rect 28586 31912 28680 31940
rect 31476 32236 31570 32264
rect 31476 32180 31495 32236
rect 31551 32180 31570 32236
rect 31476 32156 31570 32180
rect 31476 32100 31495 32156
rect 31551 32100 31570 32156
rect 31476 32076 31570 32100
rect 31476 32020 31495 32076
rect 31551 32020 31570 32076
rect 31476 31996 31570 32020
rect 31476 31940 31495 31996
rect 31551 31940 31570 31996
rect 31476 31912 31570 31940
rect 34366 32236 34460 32264
rect 34366 32180 34385 32236
rect 34441 32180 34460 32236
rect 34366 32156 34460 32180
rect 34366 32100 34385 32156
rect 34441 32100 34460 32156
rect 34366 32076 34460 32100
rect 34366 32020 34385 32076
rect 34441 32020 34460 32076
rect 34366 31996 34460 32020
rect 34366 31940 34385 31996
rect 34441 31940 34460 31996
rect 34366 31912 34460 31940
rect 37256 32236 37350 32264
rect 37256 32180 37275 32236
rect 37331 32180 37350 32236
rect 37256 32156 37350 32180
rect 37256 32100 37275 32156
rect 37331 32100 37350 32156
rect 37256 32076 37350 32100
rect 37256 32020 37275 32076
rect 37331 32020 37350 32076
rect 37256 31996 37350 32020
rect 37256 31940 37275 31996
rect 37331 31940 37350 31996
rect 37256 31912 37350 31940
rect 40146 32236 40240 32264
rect 40146 32180 40165 32236
rect 40221 32180 40240 32236
rect 40146 32156 40240 32180
rect 40146 32100 40165 32156
rect 40221 32100 40240 32156
rect 40146 32076 40240 32100
rect 40146 32020 40165 32076
rect 40221 32020 40240 32076
rect 40146 31996 40240 32020
rect 40146 31940 40165 31996
rect 40221 31940 40240 31996
rect 40146 31912 40240 31940
rect 43036 32236 43130 32264
rect 43036 32180 43055 32236
rect 43111 32180 43130 32236
rect 43036 32156 43130 32180
rect 43036 32100 43055 32156
rect 43111 32100 43130 32156
rect 43036 32076 43130 32100
rect 43036 32020 43055 32076
rect 43111 32020 43130 32076
rect 43036 31996 43130 32020
rect 43036 31940 43055 31996
rect 43111 31940 43130 31996
rect 43036 31912 43130 31940
rect 45926 32236 46020 32264
rect 45926 32180 45945 32236
rect 46001 32180 46020 32236
rect 45926 32156 46020 32180
rect 45926 32100 45945 32156
rect 46001 32100 46020 32156
rect 45926 32076 46020 32100
rect 45926 32020 45945 32076
rect 46001 32020 46020 32076
rect 45926 31996 46020 32020
rect 45926 31940 45945 31996
rect 46001 31940 46020 31996
rect 45926 31912 46020 31940
rect 48873 32236 48967 32264
rect 48873 32180 48892 32236
rect 48948 32180 48967 32236
rect 48873 32156 48967 32180
rect 48873 32100 48892 32156
rect 48948 32100 48967 32156
rect 48873 32076 48967 32100
rect 48873 32020 48892 32076
rect 48948 32020 48967 32076
rect 48873 31996 48967 32020
rect 48873 31940 48892 31996
rect 48948 31940 48967 31996
rect 48873 31912 48967 31940
rect 49722 32236 49922 32264
rect 49722 32180 49754 32236
rect 49810 32180 49834 32236
rect 49890 32180 49922 32236
rect 49722 32156 49922 32180
rect 49722 32100 49754 32156
rect 49810 32100 49834 32156
rect 49890 32100 49922 32156
rect 49722 32076 49922 32100
rect 49722 32020 49754 32076
rect 49810 32020 49834 32076
rect 49890 32020 49922 32076
rect 49722 31996 49922 32020
rect 49722 31940 49754 31996
rect 49810 31940 49834 31996
rect 49890 31940 49922 31996
rect 49722 31912 49922 31940
rect 53012 32236 53140 32264
rect 53012 32180 53048 32236
rect 53104 32180 53140 32236
rect 53012 32156 53140 32180
rect 53012 32100 53048 32156
rect 53104 32100 53140 32156
rect 53012 32076 53140 32100
rect 53012 32020 53048 32076
rect 53104 32020 53140 32076
rect 53012 31996 53140 32020
rect 53012 31940 53048 31996
rect 53104 31940 53140 31996
rect 53012 31912 53140 31940
rect 53170 32236 53298 32264
rect 53170 32180 53206 32236
rect 53262 32180 53298 32236
rect 53170 32156 53298 32180
rect 53170 32100 53206 32156
rect 53262 32100 53298 32156
rect 53170 32076 53298 32100
rect 53170 32020 53206 32076
rect 53262 32020 53298 32076
rect 53170 31996 53298 32020
rect 53170 31940 53206 31996
rect 53262 31940 53298 31996
rect 53170 31912 53298 31940
rect 53526 32236 53654 32264
rect 53526 32180 53562 32236
rect 53618 32180 53654 32236
rect 53526 32156 53654 32180
rect 53526 32100 53562 32156
rect 53618 32100 53654 32156
rect 53526 32076 53654 32100
rect 53526 32020 53562 32076
rect 53618 32020 53654 32076
rect 53526 31996 53654 32020
rect 53526 31940 53562 31996
rect 53618 31940 53654 31996
rect 53526 31912 53654 31940
rect 54844 32236 54972 32264
rect 54844 32180 54880 32236
rect 54936 32180 54972 32236
rect 54844 32156 54972 32180
rect 54844 32100 54880 32156
rect 54936 32100 54972 32156
rect 54844 32076 54972 32100
rect 54844 32020 54880 32076
rect 54936 32020 54972 32076
rect 54844 31996 54972 32020
rect 54844 31940 54880 31996
rect 54936 31940 54972 31996
rect 54844 31912 54972 31940
rect 55437 32236 55565 32264
rect 55437 32180 55473 32236
rect 55529 32180 55565 32236
rect 55437 32156 55565 32180
rect 55437 32100 55473 32156
rect 55529 32100 55565 32156
rect 55437 32076 55565 32100
rect 55437 32020 55473 32076
rect 55529 32020 55565 32076
rect 55437 31996 55565 32020
rect 55437 31940 55473 31996
rect 55529 31940 55565 31996
rect 55437 31912 55565 31940
rect 56583 32236 56711 32264
rect 56583 32180 56619 32236
rect 56675 32180 56711 32236
rect 56583 32156 56711 32180
rect 56583 32100 56619 32156
rect 56675 32100 56711 32156
rect 56583 32076 56711 32100
rect 56583 32020 56619 32076
rect 56675 32020 56711 32076
rect 56583 31996 56711 32020
rect 56583 31940 56619 31996
rect 56675 31940 56711 31996
rect 56583 31912 56711 31940
rect 58033 32236 58213 32264
rect 58033 32180 58055 32236
rect 58111 32180 58135 32236
rect 58191 32180 58213 32236
rect 58033 32156 58213 32180
rect 58033 32100 58055 32156
rect 58111 32100 58135 32156
rect 58191 32100 58213 32156
rect 58033 32076 58213 32100
rect 58033 32020 58055 32076
rect 58111 32020 58135 32076
rect 58191 32020 58213 32076
rect 58033 31996 58213 32020
rect 58033 31940 58055 31996
rect 58111 31940 58135 31996
rect 58191 31940 58213 31996
rect 58033 31912 58213 31940
rect 59256 32236 59396 32264
rect 59256 32180 59298 32236
rect 59354 32180 59396 32236
rect 59256 32156 59396 32180
rect 59256 32100 59298 32156
rect 59354 32100 59396 32156
rect 59256 32076 59396 32100
rect 59256 32020 59298 32076
rect 59354 32020 59396 32076
rect 59256 31996 59396 32020
rect 59256 31940 59298 31996
rect 59354 31940 59396 31996
rect 59256 31912 59396 31940
rect 59426 32236 59542 32264
rect 59426 32180 59456 32236
rect 59512 32180 59542 32236
rect 59426 32156 59542 32180
rect 59426 32100 59456 32156
rect 59512 32100 59542 32156
rect 59426 32076 59542 32100
rect 59426 32020 59456 32076
rect 59512 32020 59542 32076
rect 59426 31996 59542 32020
rect 59426 31940 59456 31996
rect 59512 31940 59542 31996
rect 59426 31912 59542 31940
rect 59734 32236 59850 32264
rect 59734 32180 59764 32236
rect 59820 32180 59850 32236
rect 59734 32156 59850 32180
rect 59734 32100 59764 32156
rect 59820 32100 59850 32156
rect 59734 32076 59850 32100
rect 59734 32020 59764 32076
rect 59820 32020 59850 32076
rect 59734 31996 59850 32020
rect 59734 31940 59764 31996
rect 59820 31940 59850 31996
rect 59734 31912 59850 31940
rect 59880 32236 59996 32264
rect 59880 32180 59910 32236
rect 59966 32180 59996 32236
rect 59880 32156 59996 32180
rect 59880 32100 59910 32156
rect 59966 32100 59996 32156
rect 59880 32076 59996 32100
rect 59880 32020 59910 32076
rect 59966 32020 59996 32076
rect 59880 31996 59996 32020
rect 59880 31940 59910 31996
rect 59966 31940 59996 31996
rect 59880 31912 59996 31940
rect 60026 32236 60202 32264
rect 60026 32180 60046 32236
rect 60102 32180 60126 32236
rect 60182 32180 60202 32236
rect 60026 32156 60202 32180
rect 60026 32100 60046 32156
rect 60102 32100 60126 32156
rect 60182 32100 60202 32156
rect 60026 32076 60202 32100
rect 60026 32020 60046 32076
rect 60102 32020 60126 32076
rect 60182 32020 60202 32076
rect 60026 31996 60202 32020
rect 60026 31940 60046 31996
rect 60102 31940 60126 31996
rect 60182 31940 60202 31996
rect 60026 31912 60202 31940
rect 62399 32236 62573 32264
rect 62399 32180 62418 32236
rect 62474 32180 62498 32236
rect 62554 32180 62573 32236
rect 62399 32156 62573 32180
rect 62399 32100 62418 32156
rect 62474 32100 62498 32156
rect 62554 32100 62573 32156
rect 62399 32076 62573 32100
rect 62399 32020 62418 32076
rect 62474 32020 62498 32076
rect 62554 32020 62573 32076
rect 62399 31996 62573 32020
rect 62399 31940 62418 31996
rect 62474 31940 62498 31996
rect 62554 31940 62573 31996
rect 62399 31912 62573 31940
rect 2112 24588 2216 24616
rect 2112 24532 2136 24588
rect 2192 24532 2216 24588
rect 2112 24508 2216 24532
rect 2112 24452 2136 24508
rect 2192 24452 2216 24508
rect 2112 24428 2216 24452
rect 2112 24372 2136 24428
rect 2192 24372 2216 24428
rect 2112 24348 2216 24372
rect 2112 24292 2136 24348
rect 2192 24292 2216 24348
rect 2112 24264 2216 24292
rect 5613 24588 5707 24616
rect 5613 24532 5632 24588
rect 5688 24532 5707 24588
rect 5613 24508 5707 24532
rect 5613 24452 5632 24508
rect 5688 24452 5707 24508
rect 5613 24428 5707 24452
rect 5613 24372 5632 24428
rect 5688 24372 5707 24428
rect 5613 24348 5707 24372
rect 5613 24292 5632 24348
rect 5688 24292 5707 24348
rect 5613 24264 5707 24292
rect 8503 24588 8597 24616
rect 8503 24532 8522 24588
rect 8578 24532 8597 24588
rect 8503 24508 8597 24532
rect 8503 24452 8522 24508
rect 8578 24452 8597 24508
rect 8503 24428 8597 24452
rect 8503 24372 8522 24428
rect 8578 24372 8597 24428
rect 8503 24348 8597 24372
rect 8503 24292 8522 24348
rect 8578 24292 8597 24348
rect 8503 24264 8597 24292
rect 11393 24588 11487 24616
rect 11393 24532 11412 24588
rect 11468 24532 11487 24588
rect 11393 24508 11487 24532
rect 11393 24452 11412 24508
rect 11468 24452 11487 24508
rect 11393 24428 11487 24452
rect 11393 24372 11412 24428
rect 11468 24372 11487 24428
rect 11393 24348 11487 24372
rect 11393 24292 11412 24348
rect 11468 24292 11487 24348
rect 11393 24264 11487 24292
rect 14283 24588 14377 24616
rect 14283 24532 14302 24588
rect 14358 24532 14377 24588
rect 14283 24508 14377 24532
rect 14283 24452 14302 24508
rect 14358 24452 14377 24508
rect 14283 24428 14377 24452
rect 14283 24372 14302 24428
rect 14358 24372 14377 24428
rect 14283 24348 14377 24372
rect 14283 24292 14302 24348
rect 14358 24292 14377 24348
rect 14283 24264 14377 24292
rect 17173 24588 17267 24616
rect 17173 24532 17192 24588
rect 17248 24532 17267 24588
rect 17173 24508 17267 24532
rect 17173 24452 17192 24508
rect 17248 24452 17267 24508
rect 17173 24428 17267 24452
rect 17173 24372 17192 24428
rect 17248 24372 17267 24428
rect 17173 24348 17267 24372
rect 17173 24292 17192 24348
rect 17248 24292 17267 24348
rect 17173 24264 17267 24292
rect 20063 24588 20157 24616
rect 20063 24532 20082 24588
rect 20138 24532 20157 24588
rect 20063 24508 20157 24532
rect 20063 24452 20082 24508
rect 20138 24452 20157 24508
rect 20063 24428 20157 24452
rect 20063 24372 20082 24428
rect 20138 24372 20157 24428
rect 20063 24348 20157 24372
rect 20063 24292 20082 24348
rect 20138 24292 20157 24348
rect 20063 24264 20157 24292
rect 22953 24588 23047 24616
rect 22953 24532 22972 24588
rect 23028 24532 23047 24588
rect 22953 24508 23047 24532
rect 22953 24452 22972 24508
rect 23028 24452 23047 24508
rect 22953 24428 23047 24452
rect 22953 24372 22972 24428
rect 23028 24372 23047 24428
rect 22953 24348 23047 24372
rect 22953 24292 22972 24348
rect 23028 24292 23047 24348
rect 22953 24264 23047 24292
rect 25843 24588 25937 24616
rect 25843 24532 25862 24588
rect 25918 24532 25937 24588
rect 25843 24508 25937 24532
rect 25843 24452 25862 24508
rect 25918 24452 25937 24508
rect 25843 24428 25937 24452
rect 25843 24372 25862 24428
rect 25918 24372 25937 24428
rect 25843 24348 25937 24372
rect 25843 24292 25862 24348
rect 25918 24292 25937 24348
rect 25843 24264 25937 24292
rect 28733 24588 28827 24616
rect 28733 24532 28752 24588
rect 28808 24532 28827 24588
rect 28733 24508 28827 24532
rect 28733 24452 28752 24508
rect 28808 24452 28827 24508
rect 28733 24428 28827 24452
rect 28733 24372 28752 24428
rect 28808 24372 28827 24428
rect 28733 24348 28827 24372
rect 28733 24292 28752 24348
rect 28808 24292 28827 24348
rect 28733 24264 28827 24292
rect 31623 24588 31717 24616
rect 31623 24532 31642 24588
rect 31698 24532 31717 24588
rect 31623 24508 31717 24532
rect 31623 24452 31642 24508
rect 31698 24452 31717 24508
rect 31623 24428 31717 24452
rect 31623 24372 31642 24428
rect 31698 24372 31717 24428
rect 31623 24348 31717 24372
rect 31623 24292 31642 24348
rect 31698 24292 31717 24348
rect 31623 24264 31717 24292
rect 34513 24588 34607 24616
rect 34513 24532 34532 24588
rect 34588 24532 34607 24588
rect 34513 24508 34607 24532
rect 34513 24452 34532 24508
rect 34588 24452 34607 24508
rect 34513 24428 34607 24452
rect 34513 24372 34532 24428
rect 34588 24372 34607 24428
rect 34513 24348 34607 24372
rect 34513 24292 34532 24348
rect 34588 24292 34607 24348
rect 34513 24264 34607 24292
rect 37403 24588 37497 24616
rect 37403 24532 37422 24588
rect 37478 24532 37497 24588
rect 37403 24508 37497 24532
rect 37403 24452 37422 24508
rect 37478 24452 37497 24508
rect 37403 24428 37497 24452
rect 37403 24372 37422 24428
rect 37478 24372 37497 24428
rect 37403 24348 37497 24372
rect 37403 24292 37422 24348
rect 37478 24292 37497 24348
rect 37403 24264 37497 24292
rect 40293 24588 40387 24616
rect 40293 24532 40312 24588
rect 40368 24532 40387 24588
rect 40293 24508 40387 24532
rect 40293 24452 40312 24508
rect 40368 24452 40387 24508
rect 40293 24428 40387 24452
rect 40293 24372 40312 24428
rect 40368 24372 40387 24428
rect 40293 24348 40387 24372
rect 40293 24292 40312 24348
rect 40368 24292 40387 24348
rect 40293 24264 40387 24292
rect 43183 24588 43277 24616
rect 43183 24532 43202 24588
rect 43258 24532 43277 24588
rect 43183 24508 43277 24532
rect 43183 24452 43202 24508
rect 43258 24452 43277 24508
rect 43183 24428 43277 24452
rect 43183 24372 43202 24428
rect 43258 24372 43277 24428
rect 43183 24348 43277 24372
rect 43183 24292 43202 24348
rect 43258 24292 43277 24348
rect 43183 24264 43277 24292
rect 46073 24588 46167 24616
rect 46073 24532 46092 24588
rect 46148 24532 46167 24588
rect 46073 24508 46167 24532
rect 46073 24452 46092 24508
rect 46148 24452 46167 24508
rect 46073 24428 46167 24452
rect 46073 24372 46092 24428
rect 46148 24372 46167 24428
rect 46073 24348 46167 24372
rect 46073 24292 46092 24348
rect 46148 24292 46167 24348
rect 46073 24264 46167 24292
rect 49081 24588 49175 24616
rect 49081 24532 49100 24588
rect 49156 24532 49175 24588
rect 49081 24508 49175 24532
rect 49081 24452 49100 24508
rect 49156 24452 49175 24508
rect 49081 24428 49175 24452
rect 49081 24372 49100 24428
rect 49156 24372 49175 24428
rect 49081 24348 49175 24372
rect 49081 24292 49100 24348
rect 49156 24292 49175 24348
rect 49081 24264 49175 24292
rect 52302 24588 52412 24616
rect 52302 24532 52329 24588
rect 52385 24532 52412 24588
rect 52302 24508 52412 24532
rect 52302 24452 52329 24508
rect 52385 24452 52412 24508
rect 52302 24428 52412 24452
rect 52302 24372 52329 24428
rect 52385 24372 52412 24428
rect 52302 24348 52412 24372
rect 52302 24292 52329 24348
rect 52385 24292 52412 24348
rect 52302 24264 52412 24292
rect 53694 24588 53822 24616
rect 53694 24532 53730 24588
rect 53786 24532 53822 24588
rect 53694 24508 53822 24532
rect 53694 24452 53730 24508
rect 53786 24452 53822 24508
rect 53694 24428 53822 24452
rect 53694 24372 53730 24428
rect 53786 24372 53822 24428
rect 53694 24348 53822 24372
rect 53694 24292 53730 24348
rect 53786 24292 53822 24348
rect 53694 24264 53822 24292
rect 53862 24588 53990 24616
rect 53862 24532 53898 24588
rect 53954 24532 53990 24588
rect 53862 24508 53990 24532
rect 53862 24452 53898 24508
rect 53954 24452 53990 24508
rect 53862 24428 53990 24452
rect 53862 24372 53898 24428
rect 53954 24372 53990 24428
rect 53862 24348 53990 24372
rect 53862 24292 53898 24348
rect 53954 24292 53990 24348
rect 53862 24264 53990 24292
rect 54606 24588 54734 24616
rect 54606 24532 54642 24588
rect 54698 24532 54734 24588
rect 54606 24508 54734 24532
rect 54606 24452 54642 24508
rect 54698 24452 54734 24508
rect 54606 24428 54734 24452
rect 54606 24372 54642 24428
rect 54698 24372 54734 24428
rect 54606 24348 54734 24372
rect 54606 24292 54642 24348
rect 54698 24292 54734 24348
rect 54606 24264 54734 24292
rect 55002 24588 55118 24616
rect 55002 24532 55032 24588
rect 55088 24532 55118 24588
rect 55002 24508 55118 24532
rect 55002 24452 55032 24508
rect 55088 24452 55118 24508
rect 55002 24428 55118 24452
rect 55002 24372 55032 24428
rect 55088 24372 55118 24428
rect 55002 24348 55118 24372
rect 55002 24292 55032 24348
rect 55088 24292 55118 24348
rect 55002 24264 55118 24292
rect 55712 24588 55840 24616
rect 55712 24532 55748 24588
rect 55804 24532 55840 24588
rect 55712 24508 55840 24532
rect 55712 24452 55748 24508
rect 55804 24452 55840 24508
rect 55712 24428 55840 24452
rect 55712 24372 55748 24428
rect 55804 24372 55840 24428
rect 55712 24348 55840 24372
rect 55712 24292 55748 24348
rect 55804 24292 55840 24348
rect 55712 24264 55840 24292
rect 56290 24588 56418 24616
rect 56290 24532 56326 24588
rect 56382 24532 56418 24588
rect 56290 24508 56418 24532
rect 56290 24452 56326 24508
rect 56382 24452 56418 24508
rect 56290 24428 56418 24452
rect 56290 24372 56326 24428
rect 56382 24372 56418 24428
rect 56290 24348 56418 24372
rect 56290 24292 56326 24348
rect 56382 24292 56418 24348
rect 56290 24264 56418 24292
rect 56741 24588 56857 24616
rect 56741 24532 56771 24588
rect 56827 24532 56857 24588
rect 56741 24508 56857 24532
rect 56741 24452 56771 24508
rect 56827 24452 56857 24508
rect 56741 24428 56857 24452
rect 56741 24372 56771 24428
rect 56827 24372 56857 24428
rect 56741 24348 56857 24372
rect 56741 24292 56771 24348
rect 56827 24292 56857 24348
rect 56741 24264 56857 24292
rect 57045 24588 57161 24616
rect 57045 24532 57075 24588
rect 57131 24532 57161 24588
rect 57045 24508 57161 24532
rect 57045 24452 57075 24508
rect 57131 24452 57161 24508
rect 57045 24428 57161 24452
rect 57045 24372 57075 24428
rect 57131 24372 57161 24428
rect 57045 24348 57161 24372
rect 57045 24292 57075 24348
rect 57131 24292 57161 24348
rect 57045 24264 57161 24292
rect 57887 24588 58003 24616
rect 57887 24532 57917 24588
rect 57973 24532 58003 24588
rect 57887 24508 58003 24532
rect 57887 24452 57917 24508
rect 57973 24452 58003 24508
rect 57887 24428 58003 24452
rect 57887 24372 57917 24428
rect 57973 24372 58003 24428
rect 57887 24348 58003 24372
rect 57887 24292 57917 24348
rect 57973 24292 58003 24348
rect 57887 24264 58003 24292
rect 58553 24588 58617 24616
rect 58553 24532 58557 24588
rect 58613 24532 58617 24588
rect 58553 24508 58617 24532
rect 58553 24452 58557 24508
rect 58613 24452 58617 24508
rect 58553 24428 58617 24452
rect 58553 24372 58557 24428
rect 58613 24372 58617 24428
rect 58553 24348 58617 24372
rect 58553 24292 58557 24348
rect 58613 24292 58617 24348
rect 58553 24264 58617 24292
rect 59110 24588 59226 24616
rect 59110 24532 59140 24588
rect 59196 24532 59226 24588
rect 59110 24508 59226 24532
rect 59110 24452 59140 24508
rect 59196 24452 59226 24508
rect 59110 24428 59226 24452
rect 59110 24372 59140 24428
rect 59196 24372 59226 24428
rect 59110 24348 59226 24372
rect 59110 24292 59140 24348
rect 59196 24292 59226 24348
rect 59110 24264 59226 24292
rect 60388 24588 60504 24616
rect 60388 24532 60418 24588
rect 60474 24532 60504 24588
rect 60388 24508 60504 24532
rect 60388 24452 60418 24508
rect 60474 24452 60504 24508
rect 60388 24428 60504 24452
rect 60388 24372 60418 24428
rect 60474 24372 60504 24428
rect 60388 24348 60504 24372
rect 60388 24292 60418 24348
rect 60474 24292 60504 24348
rect 60388 24264 60504 24292
rect 60546 24588 60662 24616
rect 60546 24532 60576 24588
rect 60632 24532 60662 24588
rect 60546 24508 60662 24532
rect 60546 24452 60576 24508
rect 60632 24452 60662 24508
rect 60546 24428 60662 24452
rect 60546 24372 60576 24428
rect 60632 24372 60662 24428
rect 60546 24348 60662 24372
rect 60546 24292 60576 24348
rect 60632 24292 60662 24348
rect 60546 24264 60662 24292
rect 62601 24588 62775 24616
rect 62601 24532 62620 24588
rect 62676 24532 62700 24588
rect 62756 24532 62775 24588
rect 62601 24508 62775 24532
rect 62601 24452 62620 24508
rect 62676 24452 62700 24508
rect 62756 24452 62775 24508
rect 62601 24428 62775 24452
rect 62601 24372 62620 24428
rect 62676 24372 62700 24428
rect 62756 24372 62775 24428
rect 62601 24348 62775 24372
rect 62601 24292 62620 24348
rect 62676 24292 62700 24348
rect 62756 24292 62775 24348
rect 62601 24264 62775 24292
rect 63512 22778 63540 37810
rect 63500 22772 63552 22778
rect 63500 22714 63552 22720
rect 63500 22568 63552 22574
rect 63500 22510 63552 22516
rect 2244 22236 2444 22264
rect 2244 22180 2276 22236
rect 2332 22180 2356 22236
rect 2412 22180 2444 22236
rect 2244 22156 2444 22180
rect 2244 22100 2276 22156
rect 2332 22100 2356 22156
rect 2412 22100 2444 22156
rect 2244 22076 2444 22100
rect 2244 22020 2276 22076
rect 2332 22020 2356 22076
rect 2412 22020 2444 22076
rect 2244 21996 2444 22020
rect 2244 21940 2276 21996
rect 2332 21940 2356 21996
rect 2412 21940 2444 21996
rect 2244 21912 2444 21940
rect 5466 22236 5560 22264
rect 5466 22180 5485 22236
rect 5541 22180 5560 22236
rect 5466 22156 5560 22180
rect 5466 22100 5485 22156
rect 5541 22100 5560 22156
rect 5466 22076 5560 22100
rect 5466 22020 5485 22076
rect 5541 22020 5560 22076
rect 5466 21996 5560 22020
rect 5466 21940 5485 21996
rect 5541 21940 5560 21996
rect 5466 21912 5560 21940
rect 8356 22236 8450 22264
rect 8356 22180 8375 22236
rect 8431 22180 8450 22236
rect 8356 22156 8450 22180
rect 8356 22100 8375 22156
rect 8431 22100 8450 22156
rect 8356 22076 8450 22100
rect 8356 22020 8375 22076
rect 8431 22020 8450 22076
rect 8356 21996 8450 22020
rect 8356 21940 8375 21996
rect 8431 21940 8450 21996
rect 8356 21912 8450 21940
rect 11246 22236 11340 22264
rect 11246 22180 11265 22236
rect 11321 22180 11340 22236
rect 11246 22156 11340 22180
rect 11246 22100 11265 22156
rect 11321 22100 11340 22156
rect 11246 22076 11340 22100
rect 11246 22020 11265 22076
rect 11321 22020 11340 22076
rect 11246 21996 11340 22020
rect 11246 21940 11265 21996
rect 11321 21940 11340 21996
rect 11246 21912 11340 21940
rect 14136 22236 14230 22264
rect 14136 22180 14155 22236
rect 14211 22180 14230 22236
rect 14136 22156 14230 22180
rect 14136 22100 14155 22156
rect 14211 22100 14230 22156
rect 14136 22076 14230 22100
rect 14136 22020 14155 22076
rect 14211 22020 14230 22076
rect 14136 21996 14230 22020
rect 14136 21940 14155 21996
rect 14211 21940 14230 21996
rect 14136 21912 14230 21940
rect 17026 22236 17120 22264
rect 17026 22180 17045 22236
rect 17101 22180 17120 22236
rect 17026 22156 17120 22180
rect 17026 22100 17045 22156
rect 17101 22100 17120 22156
rect 17026 22076 17120 22100
rect 17026 22020 17045 22076
rect 17101 22020 17120 22076
rect 17026 21996 17120 22020
rect 17026 21940 17045 21996
rect 17101 21940 17120 21996
rect 17026 21912 17120 21940
rect 19916 22236 20010 22264
rect 19916 22180 19935 22236
rect 19991 22180 20010 22236
rect 19916 22156 20010 22180
rect 19916 22100 19935 22156
rect 19991 22100 20010 22156
rect 19916 22076 20010 22100
rect 19916 22020 19935 22076
rect 19991 22020 20010 22076
rect 19916 21996 20010 22020
rect 19916 21940 19935 21996
rect 19991 21940 20010 21996
rect 19916 21912 20010 21940
rect 22806 22236 22900 22264
rect 22806 22180 22825 22236
rect 22881 22180 22900 22236
rect 22806 22156 22900 22180
rect 22806 22100 22825 22156
rect 22881 22100 22900 22156
rect 22806 22076 22900 22100
rect 22806 22020 22825 22076
rect 22881 22020 22900 22076
rect 22806 21996 22900 22020
rect 22806 21940 22825 21996
rect 22881 21940 22900 21996
rect 22806 21912 22900 21940
rect 25696 22236 25790 22264
rect 25696 22180 25715 22236
rect 25771 22180 25790 22236
rect 25696 22156 25790 22180
rect 25696 22100 25715 22156
rect 25771 22100 25790 22156
rect 25696 22076 25790 22100
rect 25696 22020 25715 22076
rect 25771 22020 25790 22076
rect 25696 21996 25790 22020
rect 25696 21940 25715 21996
rect 25771 21940 25790 21996
rect 25696 21912 25790 21940
rect 28586 22236 28680 22264
rect 28586 22180 28605 22236
rect 28661 22180 28680 22236
rect 28586 22156 28680 22180
rect 28586 22100 28605 22156
rect 28661 22100 28680 22156
rect 28586 22076 28680 22100
rect 28586 22020 28605 22076
rect 28661 22020 28680 22076
rect 28586 21996 28680 22020
rect 28586 21940 28605 21996
rect 28661 21940 28680 21996
rect 28586 21912 28680 21940
rect 31476 22236 31570 22264
rect 31476 22180 31495 22236
rect 31551 22180 31570 22236
rect 31476 22156 31570 22180
rect 31476 22100 31495 22156
rect 31551 22100 31570 22156
rect 31476 22076 31570 22100
rect 31476 22020 31495 22076
rect 31551 22020 31570 22076
rect 31476 21996 31570 22020
rect 31476 21940 31495 21996
rect 31551 21940 31570 21996
rect 31476 21912 31570 21940
rect 34366 22236 34460 22264
rect 34366 22180 34385 22236
rect 34441 22180 34460 22236
rect 34366 22156 34460 22180
rect 34366 22100 34385 22156
rect 34441 22100 34460 22156
rect 34366 22076 34460 22100
rect 34366 22020 34385 22076
rect 34441 22020 34460 22076
rect 34366 21996 34460 22020
rect 34366 21940 34385 21996
rect 34441 21940 34460 21996
rect 34366 21912 34460 21940
rect 37256 22236 37350 22264
rect 37256 22180 37275 22236
rect 37331 22180 37350 22236
rect 37256 22156 37350 22180
rect 37256 22100 37275 22156
rect 37331 22100 37350 22156
rect 37256 22076 37350 22100
rect 37256 22020 37275 22076
rect 37331 22020 37350 22076
rect 37256 21996 37350 22020
rect 37256 21940 37275 21996
rect 37331 21940 37350 21996
rect 37256 21912 37350 21940
rect 40146 22236 40240 22264
rect 40146 22180 40165 22236
rect 40221 22180 40240 22236
rect 40146 22156 40240 22180
rect 40146 22100 40165 22156
rect 40221 22100 40240 22156
rect 40146 22076 40240 22100
rect 40146 22020 40165 22076
rect 40221 22020 40240 22076
rect 40146 21996 40240 22020
rect 40146 21940 40165 21996
rect 40221 21940 40240 21996
rect 40146 21912 40240 21940
rect 43036 22236 43130 22264
rect 43036 22180 43055 22236
rect 43111 22180 43130 22236
rect 43036 22156 43130 22180
rect 43036 22100 43055 22156
rect 43111 22100 43130 22156
rect 43036 22076 43130 22100
rect 43036 22020 43055 22076
rect 43111 22020 43130 22076
rect 43036 21996 43130 22020
rect 43036 21940 43055 21996
rect 43111 21940 43130 21996
rect 43036 21912 43130 21940
rect 45926 22236 46020 22264
rect 45926 22180 45945 22236
rect 46001 22180 46020 22236
rect 45926 22156 46020 22180
rect 45926 22100 45945 22156
rect 46001 22100 46020 22156
rect 45926 22076 46020 22100
rect 45926 22020 45945 22076
rect 46001 22020 46020 22076
rect 45926 21996 46020 22020
rect 45926 21940 45945 21996
rect 46001 21940 46020 21996
rect 45926 21912 46020 21940
rect 48873 22236 48967 22264
rect 48873 22180 48892 22236
rect 48948 22180 48967 22236
rect 48873 22156 48967 22180
rect 48873 22100 48892 22156
rect 48948 22100 48967 22156
rect 48873 22076 48967 22100
rect 48873 22020 48892 22076
rect 48948 22020 48967 22076
rect 48873 21996 48967 22020
rect 48873 21940 48892 21996
rect 48948 21940 48967 21996
rect 48873 21912 48967 21940
rect 49722 22236 49922 22264
rect 49722 22180 49754 22236
rect 49810 22180 49834 22236
rect 49890 22180 49922 22236
rect 49722 22156 49922 22180
rect 49722 22100 49754 22156
rect 49810 22100 49834 22156
rect 49890 22100 49922 22156
rect 49722 22076 49922 22100
rect 49722 22020 49754 22076
rect 49810 22020 49834 22076
rect 49890 22020 49922 22076
rect 49722 21996 49922 22020
rect 49722 21940 49754 21996
rect 49810 21940 49834 21996
rect 49890 21940 49922 21996
rect 49722 21912 49922 21940
rect 53012 22236 53140 22264
rect 53012 22180 53048 22236
rect 53104 22180 53140 22236
rect 53012 22156 53140 22180
rect 53012 22100 53048 22156
rect 53104 22100 53140 22156
rect 53012 22076 53140 22100
rect 53012 22020 53048 22076
rect 53104 22020 53140 22076
rect 53012 21996 53140 22020
rect 53012 21940 53048 21996
rect 53104 21940 53140 21996
rect 53012 21912 53140 21940
rect 53170 22236 53298 22264
rect 53170 22180 53206 22236
rect 53262 22180 53298 22236
rect 53170 22156 53298 22180
rect 53170 22100 53206 22156
rect 53262 22100 53298 22156
rect 53170 22076 53298 22100
rect 53170 22020 53206 22076
rect 53262 22020 53298 22076
rect 53170 21996 53298 22020
rect 53170 21940 53206 21996
rect 53262 21940 53298 21996
rect 53170 21912 53298 21940
rect 53526 22236 53654 22264
rect 53526 22180 53562 22236
rect 53618 22180 53654 22236
rect 53526 22156 53654 22180
rect 53526 22100 53562 22156
rect 53618 22100 53654 22156
rect 53526 22076 53654 22100
rect 53526 22020 53562 22076
rect 53618 22020 53654 22076
rect 53526 21996 53654 22020
rect 53526 21940 53562 21996
rect 53618 21940 53654 21996
rect 53526 21912 53654 21940
rect 54844 22236 54972 22264
rect 54844 22180 54880 22236
rect 54936 22180 54972 22236
rect 54844 22156 54972 22180
rect 54844 22100 54880 22156
rect 54936 22100 54972 22156
rect 54844 22076 54972 22100
rect 54844 22020 54880 22076
rect 54936 22020 54972 22076
rect 54844 21996 54972 22020
rect 54844 21940 54880 21996
rect 54936 21940 54972 21996
rect 54844 21912 54972 21940
rect 55437 22236 55565 22264
rect 55437 22180 55473 22236
rect 55529 22180 55565 22236
rect 55437 22156 55565 22180
rect 55437 22100 55473 22156
rect 55529 22100 55565 22156
rect 55437 22076 55565 22100
rect 55437 22020 55473 22076
rect 55529 22020 55565 22076
rect 55437 21996 55565 22020
rect 55437 21940 55473 21996
rect 55529 21940 55565 21996
rect 55437 21912 55565 21940
rect 56583 22236 56711 22264
rect 56583 22180 56619 22236
rect 56675 22180 56711 22236
rect 56583 22156 56711 22180
rect 56583 22100 56619 22156
rect 56675 22100 56711 22156
rect 56583 22076 56711 22100
rect 56583 22020 56619 22076
rect 56675 22020 56711 22076
rect 56583 21996 56711 22020
rect 56583 21940 56619 21996
rect 56675 21940 56711 21996
rect 56583 21912 56711 21940
rect 58033 22236 58213 22264
rect 58033 22180 58055 22236
rect 58111 22180 58135 22236
rect 58191 22180 58213 22236
rect 58033 22156 58213 22180
rect 58033 22100 58055 22156
rect 58111 22100 58135 22156
rect 58191 22100 58213 22156
rect 58033 22076 58213 22100
rect 58033 22020 58055 22076
rect 58111 22020 58135 22076
rect 58191 22020 58213 22076
rect 58033 21996 58213 22020
rect 58033 21940 58055 21996
rect 58111 21940 58135 21996
rect 58191 21940 58213 21996
rect 58033 21912 58213 21940
rect 59256 22236 59396 22264
rect 59256 22180 59298 22236
rect 59354 22180 59396 22236
rect 59256 22156 59396 22180
rect 59256 22100 59298 22156
rect 59354 22100 59396 22156
rect 59256 22076 59396 22100
rect 59256 22020 59298 22076
rect 59354 22020 59396 22076
rect 59256 21996 59396 22020
rect 59256 21940 59298 21996
rect 59354 21940 59396 21996
rect 59256 21912 59396 21940
rect 59426 22236 59542 22264
rect 59426 22180 59456 22236
rect 59512 22180 59542 22236
rect 59426 22156 59542 22180
rect 59426 22100 59456 22156
rect 59512 22100 59542 22156
rect 59426 22076 59542 22100
rect 59426 22020 59456 22076
rect 59512 22020 59542 22076
rect 59426 21996 59542 22020
rect 59426 21940 59456 21996
rect 59512 21940 59542 21996
rect 59426 21912 59542 21940
rect 59734 22236 59850 22264
rect 59734 22180 59764 22236
rect 59820 22180 59850 22236
rect 59734 22156 59850 22180
rect 59734 22100 59764 22156
rect 59820 22100 59850 22156
rect 59734 22076 59850 22100
rect 59734 22020 59764 22076
rect 59820 22020 59850 22076
rect 59734 21996 59850 22020
rect 59734 21940 59764 21996
rect 59820 21940 59850 21996
rect 59734 21912 59850 21940
rect 59880 22236 59996 22264
rect 59880 22180 59910 22236
rect 59966 22180 59996 22236
rect 59880 22156 59996 22180
rect 59880 22100 59910 22156
rect 59966 22100 59996 22156
rect 59880 22076 59996 22100
rect 59880 22020 59910 22076
rect 59966 22020 59996 22076
rect 59880 21996 59996 22020
rect 59880 21940 59910 21996
rect 59966 21940 59996 21996
rect 59880 21912 59996 21940
rect 60026 22236 60202 22264
rect 60026 22180 60046 22236
rect 60102 22180 60126 22236
rect 60182 22180 60202 22236
rect 60026 22156 60202 22180
rect 60026 22100 60046 22156
rect 60102 22100 60126 22156
rect 60182 22100 60202 22156
rect 60026 22076 60202 22100
rect 60026 22020 60046 22076
rect 60102 22020 60126 22076
rect 60182 22020 60202 22076
rect 60026 21996 60202 22020
rect 60026 21940 60046 21996
rect 60102 21940 60126 21996
rect 60182 21940 60202 21996
rect 60026 21912 60202 21940
rect 62399 22236 62573 22264
rect 62399 22180 62418 22236
rect 62474 22180 62498 22236
rect 62554 22180 62573 22236
rect 62399 22156 62573 22180
rect 62399 22100 62418 22156
rect 62474 22100 62498 22156
rect 62554 22100 62573 22156
rect 62399 22076 62573 22100
rect 62399 22020 62418 22076
rect 62474 22020 62498 22076
rect 62554 22020 62573 22076
rect 62399 21996 62573 22020
rect 62399 21940 62418 21996
rect 62474 21940 62498 21996
rect 62554 21940 62573 21996
rect 62399 21912 62573 21940
rect 63512 21350 63540 22510
rect 63500 21344 63552 21350
rect 63500 21286 63552 21292
rect 63500 21244 63552 21250
rect 63500 21186 63552 21192
rect 2112 14588 2216 14616
rect 2112 14532 2136 14588
rect 2192 14532 2216 14588
rect 2112 14508 2216 14532
rect 2112 14452 2136 14508
rect 2192 14452 2216 14508
rect 2112 14428 2216 14452
rect 2112 14372 2136 14428
rect 2192 14372 2216 14428
rect 2112 14348 2216 14372
rect 2112 14292 2136 14348
rect 2192 14292 2216 14348
rect 2112 14264 2216 14292
rect 5613 14588 5707 14616
rect 5613 14532 5632 14588
rect 5688 14532 5707 14588
rect 5613 14508 5707 14532
rect 5613 14452 5632 14508
rect 5688 14452 5707 14508
rect 5613 14428 5707 14452
rect 5613 14372 5632 14428
rect 5688 14372 5707 14428
rect 5613 14348 5707 14372
rect 5613 14292 5632 14348
rect 5688 14292 5707 14348
rect 5613 14264 5707 14292
rect 8503 14588 8597 14616
rect 8503 14532 8522 14588
rect 8578 14532 8597 14588
rect 8503 14508 8597 14532
rect 8503 14452 8522 14508
rect 8578 14452 8597 14508
rect 8503 14428 8597 14452
rect 8503 14372 8522 14428
rect 8578 14372 8597 14428
rect 8503 14348 8597 14372
rect 8503 14292 8522 14348
rect 8578 14292 8597 14348
rect 8503 14264 8597 14292
rect 11393 14588 11487 14616
rect 11393 14532 11412 14588
rect 11468 14532 11487 14588
rect 11393 14508 11487 14532
rect 11393 14452 11412 14508
rect 11468 14452 11487 14508
rect 11393 14428 11487 14452
rect 11393 14372 11412 14428
rect 11468 14372 11487 14428
rect 11393 14348 11487 14372
rect 11393 14292 11412 14348
rect 11468 14292 11487 14348
rect 11393 14264 11487 14292
rect 14283 14588 14377 14616
rect 14283 14532 14302 14588
rect 14358 14532 14377 14588
rect 14283 14508 14377 14532
rect 14283 14452 14302 14508
rect 14358 14452 14377 14508
rect 14283 14428 14377 14452
rect 14283 14372 14302 14428
rect 14358 14372 14377 14428
rect 14283 14348 14377 14372
rect 14283 14292 14302 14348
rect 14358 14292 14377 14348
rect 14283 14264 14377 14292
rect 17173 14588 17267 14616
rect 17173 14532 17192 14588
rect 17248 14532 17267 14588
rect 17173 14508 17267 14532
rect 17173 14452 17192 14508
rect 17248 14452 17267 14508
rect 17173 14428 17267 14452
rect 17173 14372 17192 14428
rect 17248 14372 17267 14428
rect 17173 14348 17267 14372
rect 17173 14292 17192 14348
rect 17248 14292 17267 14348
rect 17173 14264 17267 14292
rect 20063 14588 20157 14616
rect 20063 14532 20082 14588
rect 20138 14532 20157 14588
rect 20063 14508 20157 14532
rect 20063 14452 20082 14508
rect 20138 14452 20157 14508
rect 20063 14428 20157 14452
rect 20063 14372 20082 14428
rect 20138 14372 20157 14428
rect 20063 14348 20157 14372
rect 20063 14292 20082 14348
rect 20138 14292 20157 14348
rect 20063 14264 20157 14292
rect 22953 14588 23047 14616
rect 22953 14532 22972 14588
rect 23028 14532 23047 14588
rect 22953 14508 23047 14532
rect 22953 14452 22972 14508
rect 23028 14452 23047 14508
rect 22953 14428 23047 14452
rect 22953 14372 22972 14428
rect 23028 14372 23047 14428
rect 22953 14348 23047 14372
rect 22953 14292 22972 14348
rect 23028 14292 23047 14348
rect 22953 14264 23047 14292
rect 25843 14588 25937 14616
rect 25843 14532 25862 14588
rect 25918 14532 25937 14588
rect 25843 14508 25937 14532
rect 25843 14452 25862 14508
rect 25918 14452 25937 14508
rect 25843 14428 25937 14452
rect 25843 14372 25862 14428
rect 25918 14372 25937 14428
rect 25843 14348 25937 14372
rect 25843 14292 25862 14348
rect 25918 14292 25937 14348
rect 25843 14264 25937 14292
rect 28733 14588 28827 14616
rect 28733 14532 28752 14588
rect 28808 14532 28827 14588
rect 28733 14508 28827 14532
rect 28733 14452 28752 14508
rect 28808 14452 28827 14508
rect 28733 14428 28827 14452
rect 28733 14372 28752 14428
rect 28808 14372 28827 14428
rect 28733 14348 28827 14372
rect 28733 14292 28752 14348
rect 28808 14292 28827 14348
rect 28733 14264 28827 14292
rect 31623 14588 31717 14616
rect 31623 14532 31642 14588
rect 31698 14532 31717 14588
rect 31623 14508 31717 14532
rect 31623 14452 31642 14508
rect 31698 14452 31717 14508
rect 31623 14428 31717 14452
rect 31623 14372 31642 14428
rect 31698 14372 31717 14428
rect 31623 14348 31717 14372
rect 31623 14292 31642 14348
rect 31698 14292 31717 14348
rect 31623 14264 31717 14292
rect 34513 14588 34607 14616
rect 34513 14532 34532 14588
rect 34588 14532 34607 14588
rect 34513 14508 34607 14532
rect 34513 14452 34532 14508
rect 34588 14452 34607 14508
rect 34513 14428 34607 14452
rect 34513 14372 34532 14428
rect 34588 14372 34607 14428
rect 34513 14348 34607 14372
rect 34513 14292 34532 14348
rect 34588 14292 34607 14348
rect 34513 14264 34607 14292
rect 37403 14588 37497 14616
rect 37403 14532 37422 14588
rect 37478 14532 37497 14588
rect 37403 14508 37497 14532
rect 37403 14452 37422 14508
rect 37478 14452 37497 14508
rect 37403 14428 37497 14452
rect 37403 14372 37422 14428
rect 37478 14372 37497 14428
rect 37403 14348 37497 14372
rect 37403 14292 37422 14348
rect 37478 14292 37497 14348
rect 37403 14264 37497 14292
rect 40293 14588 40387 14616
rect 40293 14532 40312 14588
rect 40368 14532 40387 14588
rect 40293 14508 40387 14532
rect 40293 14452 40312 14508
rect 40368 14452 40387 14508
rect 40293 14428 40387 14452
rect 40293 14372 40312 14428
rect 40368 14372 40387 14428
rect 40293 14348 40387 14372
rect 40293 14292 40312 14348
rect 40368 14292 40387 14348
rect 40293 14264 40387 14292
rect 43183 14588 43277 14616
rect 43183 14532 43202 14588
rect 43258 14532 43277 14588
rect 43183 14508 43277 14532
rect 43183 14452 43202 14508
rect 43258 14452 43277 14508
rect 43183 14428 43277 14452
rect 43183 14372 43202 14428
rect 43258 14372 43277 14428
rect 43183 14348 43277 14372
rect 43183 14292 43202 14348
rect 43258 14292 43277 14348
rect 43183 14264 43277 14292
rect 46073 14588 46167 14616
rect 46073 14532 46092 14588
rect 46148 14532 46167 14588
rect 46073 14508 46167 14532
rect 46073 14452 46092 14508
rect 46148 14452 46167 14508
rect 46073 14428 46167 14452
rect 46073 14372 46092 14428
rect 46148 14372 46167 14428
rect 46073 14348 46167 14372
rect 46073 14292 46092 14348
rect 46148 14292 46167 14348
rect 46073 14264 46167 14292
rect 49081 14588 49175 14616
rect 49081 14532 49100 14588
rect 49156 14532 49175 14588
rect 49081 14508 49175 14532
rect 49081 14452 49100 14508
rect 49156 14452 49175 14508
rect 49081 14428 49175 14452
rect 49081 14372 49100 14428
rect 49156 14372 49175 14428
rect 49081 14348 49175 14372
rect 49081 14292 49100 14348
rect 49156 14292 49175 14348
rect 49081 14264 49175 14292
rect 52302 14588 52412 14616
rect 52302 14532 52329 14588
rect 52385 14532 52412 14588
rect 52302 14508 52412 14532
rect 52302 14452 52329 14508
rect 52385 14452 52412 14508
rect 52302 14428 52412 14452
rect 52302 14372 52329 14428
rect 52385 14372 52412 14428
rect 52302 14348 52412 14372
rect 52302 14292 52329 14348
rect 52385 14292 52412 14348
rect 52302 14264 52412 14292
rect 53694 14588 53822 14616
rect 53694 14532 53730 14588
rect 53786 14532 53822 14588
rect 53694 14508 53822 14532
rect 53694 14452 53730 14508
rect 53786 14452 53822 14508
rect 53694 14428 53822 14452
rect 53694 14372 53730 14428
rect 53786 14372 53822 14428
rect 53694 14348 53822 14372
rect 53694 14292 53730 14348
rect 53786 14292 53822 14348
rect 53694 14264 53822 14292
rect 53862 14588 53990 14616
rect 53862 14532 53898 14588
rect 53954 14532 53990 14588
rect 53862 14508 53990 14532
rect 53862 14452 53898 14508
rect 53954 14452 53990 14508
rect 53862 14428 53990 14452
rect 53862 14372 53898 14428
rect 53954 14372 53990 14428
rect 53862 14348 53990 14372
rect 53862 14292 53898 14348
rect 53954 14292 53990 14348
rect 53862 14264 53990 14292
rect 54606 14588 54734 14616
rect 54606 14532 54642 14588
rect 54698 14532 54734 14588
rect 54606 14508 54734 14532
rect 54606 14452 54642 14508
rect 54698 14452 54734 14508
rect 54606 14428 54734 14452
rect 54606 14372 54642 14428
rect 54698 14372 54734 14428
rect 54606 14348 54734 14372
rect 54606 14292 54642 14348
rect 54698 14292 54734 14348
rect 54606 14264 54734 14292
rect 55002 14588 55118 14616
rect 55002 14532 55032 14588
rect 55088 14532 55118 14588
rect 55002 14508 55118 14532
rect 55002 14452 55032 14508
rect 55088 14452 55118 14508
rect 55002 14428 55118 14452
rect 55002 14372 55032 14428
rect 55088 14372 55118 14428
rect 55002 14348 55118 14372
rect 55002 14292 55032 14348
rect 55088 14292 55118 14348
rect 55002 14264 55118 14292
rect 55712 14588 55840 14616
rect 55712 14532 55748 14588
rect 55804 14532 55840 14588
rect 55712 14508 55840 14532
rect 55712 14452 55748 14508
rect 55804 14452 55840 14508
rect 55712 14428 55840 14452
rect 55712 14372 55748 14428
rect 55804 14372 55840 14428
rect 55712 14348 55840 14372
rect 55712 14292 55748 14348
rect 55804 14292 55840 14348
rect 55712 14264 55840 14292
rect 56290 14588 56418 14616
rect 56290 14532 56326 14588
rect 56382 14532 56418 14588
rect 56290 14508 56418 14532
rect 56290 14452 56326 14508
rect 56382 14452 56418 14508
rect 56290 14428 56418 14452
rect 56290 14372 56326 14428
rect 56382 14372 56418 14428
rect 56290 14348 56418 14372
rect 56290 14292 56326 14348
rect 56382 14292 56418 14348
rect 56290 14264 56418 14292
rect 56741 14588 56857 14616
rect 56741 14532 56771 14588
rect 56827 14532 56857 14588
rect 56741 14508 56857 14532
rect 56741 14452 56771 14508
rect 56827 14452 56857 14508
rect 56741 14428 56857 14452
rect 56741 14372 56771 14428
rect 56827 14372 56857 14428
rect 56741 14348 56857 14372
rect 56741 14292 56771 14348
rect 56827 14292 56857 14348
rect 56741 14264 56857 14292
rect 57045 14588 57161 14616
rect 57045 14532 57075 14588
rect 57131 14532 57161 14588
rect 57045 14508 57161 14532
rect 57045 14452 57075 14508
rect 57131 14452 57161 14508
rect 57045 14428 57161 14452
rect 57045 14372 57075 14428
rect 57131 14372 57161 14428
rect 57045 14348 57161 14372
rect 57045 14292 57075 14348
rect 57131 14292 57161 14348
rect 57045 14264 57161 14292
rect 57887 14588 58003 14616
rect 57887 14532 57917 14588
rect 57973 14532 58003 14588
rect 57887 14508 58003 14532
rect 57887 14452 57917 14508
rect 57973 14452 58003 14508
rect 57887 14428 58003 14452
rect 57887 14372 57917 14428
rect 57973 14372 58003 14428
rect 57887 14348 58003 14372
rect 57887 14292 57917 14348
rect 57973 14292 58003 14348
rect 57887 14264 58003 14292
rect 58553 14588 58617 14616
rect 58553 14532 58557 14588
rect 58613 14532 58617 14588
rect 58553 14508 58617 14532
rect 58553 14452 58557 14508
rect 58613 14452 58617 14508
rect 58553 14428 58617 14452
rect 58553 14372 58557 14428
rect 58613 14372 58617 14428
rect 58553 14348 58617 14372
rect 58553 14292 58557 14348
rect 58613 14292 58617 14348
rect 58553 14264 58617 14292
rect 59110 14588 59226 14616
rect 59110 14532 59140 14588
rect 59196 14532 59226 14588
rect 59110 14508 59226 14532
rect 59110 14452 59140 14508
rect 59196 14452 59226 14508
rect 59110 14428 59226 14452
rect 59110 14372 59140 14428
rect 59196 14372 59226 14428
rect 59110 14348 59226 14372
rect 59110 14292 59140 14348
rect 59196 14292 59226 14348
rect 59110 14264 59226 14292
rect 60388 14588 60504 14616
rect 60388 14532 60418 14588
rect 60474 14532 60504 14588
rect 60388 14508 60504 14532
rect 60388 14452 60418 14508
rect 60474 14452 60504 14508
rect 60388 14428 60504 14452
rect 60388 14372 60418 14428
rect 60474 14372 60504 14428
rect 60388 14348 60504 14372
rect 60388 14292 60418 14348
rect 60474 14292 60504 14348
rect 60388 14264 60504 14292
rect 60546 14588 60662 14616
rect 60546 14532 60576 14588
rect 60632 14532 60662 14588
rect 60546 14508 60662 14532
rect 60546 14452 60576 14508
rect 60632 14452 60662 14508
rect 60546 14428 60662 14452
rect 60546 14372 60576 14428
rect 60632 14372 60662 14428
rect 60546 14348 60662 14372
rect 60546 14292 60576 14348
rect 60632 14292 60662 14348
rect 60546 14264 60662 14292
rect 62601 14588 62775 14616
rect 62601 14532 62620 14588
rect 62676 14532 62700 14588
rect 62756 14532 62775 14588
rect 62601 14508 62775 14532
rect 62601 14452 62620 14508
rect 62676 14452 62700 14508
rect 62756 14452 62775 14508
rect 62601 14428 62775 14452
rect 62601 14372 62620 14428
rect 62676 14372 62700 14428
rect 62756 14372 62775 14428
rect 62601 14348 62775 14372
rect 62601 14292 62620 14348
rect 62676 14292 62700 14348
rect 62756 14292 62775 14348
rect 62601 14264 62775 14292
rect 2244 12236 2444 12264
rect 2244 12180 2276 12236
rect 2332 12180 2356 12236
rect 2412 12180 2444 12236
rect 2244 12156 2444 12180
rect 2244 12100 2276 12156
rect 2332 12100 2356 12156
rect 2412 12100 2444 12156
rect 2244 12076 2444 12100
rect 2244 12020 2276 12076
rect 2332 12020 2356 12076
rect 2412 12020 2444 12076
rect 2244 11996 2444 12020
rect 2244 11940 2276 11996
rect 2332 11940 2356 11996
rect 2412 11940 2444 11996
rect 2244 11912 2444 11940
rect 5466 12236 5560 12264
rect 5466 12180 5485 12236
rect 5541 12180 5560 12236
rect 5466 12156 5560 12180
rect 5466 12100 5485 12156
rect 5541 12100 5560 12156
rect 5466 12076 5560 12100
rect 5466 12020 5485 12076
rect 5541 12020 5560 12076
rect 5466 11996 5560 12020
rect 5466 11940 5485 11996
rect 5541 11940 5560 11996
rect 5466 11912 5560 11940
rect 8356 12236 8450 12264
rect 8356 12180 8375 12236
rect 8431 12180 8450 12236
rect 8356 12156 8450 12180
rect 8356 12100 8375 12156
rect 8431 12100 8450 12156
rect 8356 12076 8450 12100
rect 8356 12020 8375 12076
rect 8431 12020 8450 12076
rect 8356 11996 8450 12020
rect 8356 11940 8375 11996
rect 8431 11940 8450 11996
rect 8356 11912 8450 11940
rect 11246 12236 11340 12264
rect 11246 12180 11265 12236
rect 11321 12180 11340 12236
rect 11246 12156 11340 12180
rect 11246 12100 11265 12156
rect 11321 12100 11340 12156
rect 11246 12076 11340 12100
rect 11246 12020 11265 12076
rect 11321 12020 11340 12076
rect 11246 11996 11340 12020
rect 11246 11940 11265 11996
rect 11321 11940 11340 11996
rect 11246 11912 11340 11940
rect 14136 12236 14230 12264
rect 14136 12180 14155 12236
rect 14211 12180 14230 12236
rect 14136 12156 14230 12180
rect 14136 12100 14155 12156
rect 14211 12100 14230 12156
rect 14136 12076 14230 12100
rect 14136 12020 14155 12076
rect 14211 12020 14230 12076
rect 14136 11996 14230 12020
rect 14136 11940 14155 11996
rect 14211 11940 14230 11996
rect 14136 11912 14230 11940
rect 17026 12236 17120 12264
rect 17026 12180 17045 12236
rect 17101 12180 17120 12236
rect 17026 12156 17120 12180
rect 17026 12100 17045 12156
rect 17101 12100 17120 12156
rect 17026 12076 17120 12100
rect 17026 12020 17045 12076
rect 17101 12020 17120 12076
rect 17026 11996 17120 12020
rect 17026 11940 17045 11996
rect 17101 11940 17120 11996
rect 17026 11912 17120 11940
rect 19916 12236 20010 12264
rect 19916 12180 19935 12236
rect 19991 12180 20010 12236
rect 19916 12156 20010 12180
rect 19916 12100 19935 12156
rect 19991 12100 20010 12156
rect 19916 12076 20010 12100
rect 19916 12020 19935 12076
rect 19991 12020 20010 12076
rect 19916 11996 20010 12020
rect 19916 11940 19935 11996
rect 19991 11940 20010 11996
rect 19916 11912 20010 11940
rect 22806 12236 22900 12264
rect 22806 12180 22825 12236
rect 22881 12180 22900 12236
rect 22806 12156 22900 12180
rect 22806 12100 22825 12156
rect 22881 12100 22900 12156
rect 22806 12076 22900 12100
rect 22806 12020 22825 12076
rect 22881 12020 22900 12076
rect 22806 11996 22900 12020
rect 22806 11940 22825 11996
rect 22881 11940 22900 11996
rect 22806 11912 22900 11940
rect 25696 12236 25790 12264
rect 25696 12180 25715 12236
rect 25771 12180 25790 12236
rect 25696 12156 25790 12180
rect 25696 12100 25715 12156
rect 25771 12100 25790 12156
rect 25696 12076 25790 12100
rect 25696 12020 25715 12076
rect 25771 12020 25790 12076
rect 25696 11996 25790 12020
rect 25696 11940 25715 11996
rect 25771 11940 25790 11996
rect 25696 11912 25790 11940
rect 28586 12236 28680 12264
rect 28586 12180 28605 12236
rect 28661 12180 28680 12236
rect 28586 12156 28680 12180
rect 28586 12100 28605 12156
rect 28661 12100 28680 12156
rect 28586 12076 28680 12100
rect 28586 12020 28605 12076
rect 28661 12020 28680 12076
rect 28586 11996 28680 12020
rect 28586 11940 28605 11996
rect 28661 11940 28680 11996
rect 28586 11912 28680 11940
rect 31476 12236 31570 12264
rect 31476 12180 31495 12236
rect 31551 12180 31570 12236
rect 31476 12156 31570 12180
rect 31476 12100 31495 12156
rect 31551 12100 31570 12156
rect 31476 12076 31570 12100
rect 31476 12020 31495 12076
rect 31551 12020 31570 12076
rect 31476 11996 31570 12020
rect 31476 11940 31495 11996
rect 31551 11940 31570 11996
rect 31476 11912 31570 11940
rect 34366 12236 34460 12264
rect 34366 12180 34385 12236
rect 34441 12180 34460 12236
rect 34366 12156 34460 12180
rect 34366 12100 34385 12156
rect 34441 12100 34460 12156
rect 34366 12076 34460 12100
rect 34366 12020 34385 12076
rect 34441 12020 34460 12076
rect 34366 11996 34460 12020
rect 34366 11940 34385 11996
rect 34441 11940 34460 11996
rect 34366 11912 34460 11940
rect 37256 12236 37350 12264
rect 37256 12180 37275 12236
rect 37331 12180 37350 12236
rect 37256 12156 37350 12180
rect 37256 12100 37275 12156
rect 37331 12100 37350 12156
rect 37256 12076 37350 12100
rect 37256 12020 37275 12076
rect 37331 12020 37350 12076
rect 37256 11996 37350 12020
rect 37256 11940 37275 11996
rect 37331 11940 37350 11996
rect 37256 11912 37350 11940
rect 40146 12236 40240 12264
rect 40146 12180 40165 12236
rect 40221 12180 40240 12236
rect 40146 12156 40240 12180
rect 40146 12100 40165 12156
rect 40221 12100 40240 12156
rect 40146 12076 40240 12100
rect 40146 12020 40165 12076
rect 40221 12020 40240 12076
rect 40146 11996 40240 12020
rect 40146 11940 40165 11996
rect 40221 11940 40240 11996
rect 40146 11912 40240 11940
rect 43036 12236 43130 12264
rect 43036 12180 43055 12236
rect 43111 12180 43130 12236
rect 43036 12156 43130 12180
rect 43036 12100 43055 12156
rect 43111 12100 43130 12156
rect 43036 12076 43130 12100
rect 43036 12020 43055 12076
rect 43111 12020 43130 12076
rect 43036 11996 43130 12020
rect 43036 11940 43055 11996
rect 43111 11940 43130 11996
rect 43036 11912 43130 11940
rect 45926 12236 46020 12264
rect 45926 12180 45945 12236
rect 46001 12180 46020 12236
rect 45926 12156 46020 12180
rect 45926 12100 45945 12156
rect 46001 12100 46020 12156
rect 45926 12076 46020 12100
rect 45926 12020 45945 12076
rect 46001 12020 46020 12076
rect 45926 11996 46020 12020
rect 45926 11940 45945 11996
rect 46001 11940 46020 11996
rect 45926 11912 46020 11940
rect 48873 12236 48967 12264
rect 48873 12180 48892 12236
rect 48948 12180 48967 12236
rect 48873 12156 48967 12180
rect 48873 12100 48892 12156
rect 48948 12100 48967 12156
rect 48873 12076 48967 12100
rect 48873 12020 48892 12076
rect 48948 12020 48967 12076
rect 48873 11996 48967 12020
rect 48873 11940 48892 11996
rect 48948 11940 48967 11996
rect 48873 11912 48967 11940
rect 49722 12236 49922 12264
rect 49722 12180 49754 12236
rect 49810 12180 49834 12236
rect 49890 12180 49922 12236
rect 49722 12156 49922 12180
rect 49722 12100 49754 12156
rect 49810 12100 49834 12156
rect 49890 12100 49922 12156
rect 49722 12076 49922 12100
rect 49722 12020 49754 12076
rect 49810 12020 49834 12076
rect 49890 12020 49922 12076
rect 49722 11996 49922 12020
rect 49722 11940 49754 11996
rect 49810 11940 49834 11996
rect 49890 11940 49922 11996
rect 49722 11912 49922 11940
rect 53012 12236 53140 12264
rect 53012 12180 53048 12236
rect 53104 12180 53140 12236
rect 53012 12156 53140 12180
rect 53012 12100 53048 12156
rect 53104 12100 53140 12156
rect 53012 12076 53140 12100
rect 53012 12020 53048 12076
rect 53104 12020 53140 12076
rect 53012 11996 53140 12020
rect 53012 11940 53048 11996
rect 53104 11940 53140 11996
rect 53012 11912 53140 11940
rect 53170 12236 53298 12264
rect 53170 12180 53206 12236
rect 53262 12180 53298 12236
rect 53170 12156 53298 12180
rect 53170 12100 53206 12156
rect 53262 12100 53298 12156
rect 53170 12076 53298 12100
rect 53170 12020 53206 12076
rect 53262 12020 53298 12076
rect 53170 11996 53298 12020
rect 53170 11940 53206 11996
rect 53262 11940 53298 11996
rect 53170 11912 53298 11940
rect 53526 12236 53654 12264
rect 53526 12180 53562 12236
rect 53618 12180 53654 12236
rect 53526 12156 53654 12180
rect 53526 12100 53562 12156
rect 53618 12100 53654 12156
rect 53526 12076 53654 12100
rect 53526 12020 53562 12076
rect 53618 12020 53654 12076
rect 53526 11996 53654 12020
rect 53526 11940 53562 11996
rect 53618 11940 53654 11996
rect 53526 11912 53654 11940
rect 54844 12236 54972 12264
rect 54844 12180 54880 12236
rect 54936 12180 54972 12236
rect 54844 12156 54972 12180
rect 54844 12100 54880 12156
rect 54936 12100 54972 12156
rect 54844 12076 54972 12100
rect 54844 12020 54880 12076
rect 54936 12020 54972 12076
rect 54844 11996 54972 12020
rect 54844 11940 54880 11996
rect 54936 11940 54972 11996
rect 54844 11912 54972 11940
rect 55437 12236 55565 12264
rect 55437 12180 55473 12236
rect 55529 12180 55565 12236
rect 55437 12156 55565 12180
rect 55437 12100 55473 12156
rect 55529 12100 55565 12156
rect 55437 12076 55565 12100
rect 55437 12020 55473 12076
rect 55529 12020 55565 12076
rect 55437 11996 55565 12020
rect 55437 11940 55473 11996
rect 55529 11940 55565 11996
rect 55437 11912 55565 11940
rect 56583 12236 56711 12264
rect 56583 12180 56619 12236
rect 56675 12180 56711 12236
rect 56583 12156 56711 12180
rect 56583 12100 56619 12156
rect 56675 12100 56711 12156
rect 56583 12076 56711 12100
rect 56583 12020 56619 12076
rect 56675 12020 56711 12076
rect 56583 11996 56711 12020
rect 56583 11940 56619 11996
rect 56675 11940 56711 11996
rect 56583 11912 56711 11940
rect 58033 12236 58213 12264
rect 58033 12180 58055 12236
rect 58111 12180 58135 12236
rect 58191 12180 58213 12236
rect 58033 12156 58213 12180
rect 58033 12100 58055 12156
rect 58111 12100 58135 12156
rect 58191 12100 58213 12156
rect 58033 12076 58213 12100
rect 58033 12020 58055 12076
rect 58111 12020 58135 12076
rect 58191 12020 58213 12076
rect 58033 11996 58213 12020
rect 58033 11940 58055 11996
rect 58111 11940 58135 11996
rect 58191 11940 58213 11996
rect 58033 11912 58213 11940
rect 59256 12236 59396 12264
rect 59256 12180 59298 12236
rect 59354 12180 59396 12236
rect 59256 12156 59396 12180
rect 59256 12100 59298 12156
rect 59354 12100 59396 12156
rect 59256 12076 59396 12100
rect 59256 12020 59298 12076
rect 59354 12020 59396 12076
rect 59256 11996 59396 12020
rect 59256 11940 59298 11996
rect 59354 11940 59396 11996
rect 59256 11912 59396 11940
rect 59426 12236 59542 12264
rect 59426 12180 59456 12236
rect 59512 12180 59542 12236
rect 59426 12156 59542 12180
rect 59426 12100 59456 12156
rect 59512 12100 59542 12156
rect 59426 12076 59542 12100
rect 59426 12020 59456 12076
rect 59512 12020 59542 12076
rect 59426 11996 59542 12020
rect 59426 11940 59456 11996
rect 59512 11940 59542 11996
rect 59426 11912 59542 11940
rect 59734 12236 59850 12264
rect 59734 12180 59764 12236
rect 59820 12180 59850 12236
rect 59734 12156 59850 12180
rect 59734 12100 59764 12156
rect 59820 12100 59850 12156
rect 59734 12076 59850 12100
rect 59734 12020 59764 12076
rect 59820 12020 59850 12076
rect 59734 11996 59850 12020
rect 59734 11940 59764 11996
rect 59820 11940 59850 11996
rect 59734 11912 59850 11940
rect 59880 12236 59996 12264
rect 59880 12180 59910 12236
rect 59966 12180 59996 12236
rect 59880 12156 59996 12180
rect 59880 12100 59910 12156
rect 59966 12100 59996 12156
rect 59880 12076 59996 12100
rect 59880 12020 59910 12076
rect 59966 12020 59996 12076
rect 59880 11996 59996 12020
rect 59880 11940 59910 11996
rect 59966 11940 59996 11996
rect 59880 11912 59996 11940
rect 60026 12236 60202 12264
rect 60026 12180 60046 12236
rect 60102 12180 60126 12236
rect 60182 12180 60202 12236
rect 60026 12156 60202 12180
rect 60026 12100 60046 12156
rect 60102 12100 60126 12156
rect 60182 12100 60202 12156
rect 60026 12076 60202 12100
rect 60026 12020 60046 12076
rect 60102 12020 60126 12076
rect 60182 12020 60202 12076
rect 60026 11996 60202 12020
rect 60026 11940 60046 11996
rect 60102 11940 60126 11996
rect 60182 11940 60202 11996
rect 60026 11912 60202 11940
rect 62399 12236 62573 12264
rect 62399 12180 62418 12236
rect 62474 12180 62498 12236
rect 62554 12180 62573 12236
rect 62399 12156 62573 12180
rect 62399 12100 62418 12156
rect 62474 12100 62498 12156
rect 62554 12100 62573 12156
rect 62399 12076 62573 12100
rect 62399 12020 62418 12076
rect 62474 12020 62498 12076
rect 62554 12020 62573 12076
rect 62399 11996 62573 12020
rect 62399 11940 62418 11996
rect 62474 11940 62498 11996
rect 62554 11940 62573 11996
rect 62399 11912 62573 11940
rect 63512 10248 63540 21186
rect 63604 15881 63632 64670
rect 63696 44742 63724 76094
rect 63868 74588 63920 74594
rect 63868 74530 63920 74536
rect 63776 69624 63828 69630
rect 63776 69566 63828 69572
rect 63788 64734 63816 69566
rect 63776 64728 63828 64734
rect 63776 64670 63828 64676
rect 63776 64320 63828 64326
rect 63776 64262 63828 64268
rect 63788 62150 63816 64262
rect 63776 62144 63828 62150
rect 63776 62086 63828 62092
rect 63788 59974 63816 62086
rect 63776 59968 63828 59974
rect 63776 59910 63828 59916
rect 63788 58002 63816 59910
rect 63776 57996 63828 58002
rect 63776 57938 63828 57944
rect 63788 55622 63816 57938
rect 63776 55616 63828 55622
rect 63776 55558 63828 55564
rect 63788 53582 63816 55558
rect 63776 53576 63828 53582
rect 63776 53518 63828 53524
rect 63788 51542 63816 53518
rect 63776 51536 63828 51542
rect 63776 51478 63828 51484
rect 63684 44736 63736 44742
rect 63684 44678 63736 44684
rect 63684 44600 63736 44606
rect 63684 44542 63736 44548
rect 63696 37874 63724 44542
rect 63776 42832 63828 42838
rect 63776 42774 63828 42780
rect 63684 37868 63736 37874
rect 63684 37810 63736 37816
rect 63684 37392 63736 37398
rect 63684 37334 63736 37340
rect 63696 35222 63724 37334
rect 63684 35216 63736 35222
rect 63684 35158 63736 35164
rect 63696 33182 63724 35158
rect 63684 33176 63736 33182
rect 63684 33118 63736 33124
rect 63696 31618 63724 33118
rect 63684 31612 63736 31618
rect 63684 31554 63736 31560
rect 63684 31476 63736 31482
rect 63684 31418 63736 31424
rect 63696 23322 63724 31418
rect 63684 23316 63736 23322
rect 63684 23258 63736 23264
rect 63684 23112 63736 23118
rect 63684 23054 63736 23060
rect 63696 18193 63724 23054
rect 63682 18184 63738 18193
rect 63682 18119 63738 18128
rect 63684 18080 63736 18086
rect 63684 18022 63736 18028
rect 63590 15872 63646 15881
rect 63590 15807 63646 15816
rect 63696 15722 63724 18022
rect 63604 15694 63724 15722
rect 63604 15638 63632 15694
rect 63592 15632 63644 15638
rect 63592 15574 63644 15580
rect 63604 13734 63632 15574
rect 63592 13728 63644 13734
rect 63592 13670 63644 13676
rect 63604 11558 63632 13670
rect 63684 12436 63736 12442
rect 63684 12378 63736 12384
rect 63592 11552 63644 11558
rect 63590 11520 63592 11529
rect 63644 11520 63646 11529
rect 63590 11455 63646 11464
rect 63590 10568 63646 10577
rect 63590 10503 63646 10512
rect 63604 10350 63632 10503
rect 63592 10344 63644 10350
rect 63592 10286 63644 10292
rect 63512 10220 63632 10248
rect 63500 10056 63552 10062
rect 63498 10024 63500 10033
rect 63552 10024 63554 10033
rect 63498 9959 63554 9968
rect 63498 9888 63554 9897
rect 63498 9823 63554 9832
rect 50712 7880 50764 7886
rect 59288 7857 59316 8024
rect 50712 7822 50764 7828
rect 59274 7848 59330 7857
rect 35992 7744 36044 7750
rect 35992 7686 36044 7692
rect 32956 7608 33008 7614
rect 32956 7550 33008 7556
rect 30472 6520 30524 6526
rect 30472 6462 30524 6468
rect 30288 6452 30340 6458
rect 30288 6394 30340 6400
rect 1836 4922 2188 5944
rect 1836 4870 1858 4922
rect 1910 4870 1922 4922
rect 1974 4870 1986 4922
rect 2038 4870 2050 4922
rect 2102 4870 2114 4922
rect 2166 4870 2188 4922
rect 1836 3834 2188 4870
rect 1836 3782 1858 3834
rect 1910 3782 1922 3834
rect 1974 3782 1986 3834
rect 2038 3782 2050 3834
rect 2102 3782 2114 3834
rect 2166 3782 2188 3834
rect 1836 2746 2188 3782
rect 1836 2694 1858 2746
rect 1910 2694 1922 2746
rect 1974 2694 1986 2746
rect 2038 2694 2050 2746
rect 2102 2694 2114 2746
rect 2166 2694 2188 2746
rect 1836 2236 2188 2694
rect 1836 2180 1864 2236
rect 1920 2180 1944 2236
rect 2000 2180 2024 2236
rect 2080 2180 2104 2236
rect 2160 2180 2188 2236
rect 1836 2156 2188 2180
rect 1836 2100 1864 2156
rect 1920 2100 1944 2156
rect 2000 2100 2024 2156
rect 2080 2100 2104 2156
rect 2160 2100 2188 2156
rect 1836 2076 2188 2100
rect 1836 2020 1864 2076
rect 1920 2020 1944 2076
rect 2000 2020 2024 2076
rect 2080 2020 2104 2076
rect 2160 2020 2188 2076
rect 1836 1996 2188 2020
rect 1836 1940 1864 1996
rect 1920 1940 1944 1996
rect 2000 1940 2024 1996
rect 2080 1940 2104 1996
rect 2160 1940 2188 1996
rect 1836 1658 2188 1940
rect 1836 1606 1858 1658
rect 1910 1606 1922 1658
rect 1974 1606 1986 1658
rect 2038 1606 2050 1658
rect 2102 1606 2114 1658
rect 2166 1606 2188 1658
rect 1836 1040 2188 1606
rect 4188 5466 4540 5972
rect 4188 5414 4210 5466
rect 4262 5414 4274 5466
rect 4326 5414 4338 5466
rect 4390 5414 4402 5466
rect 4454 5414 4466 5466
rect 4518 5414 4540 5466
rect 4188 4588 4540 5414
rect 4188 4532 4216 4588
rect 4272 4532 4296 4588
rect 4352 4532 4376 4588
rect 4432 4532 4456 4588
rect 4512 4532 4540 4588
rect 4188 4508 4540 4532
rect 4188 4452 4216 4508
rect 4272 4452 4296 4508
rect 4352 4452 4376 4508
rect 4432 4452 4456 4508
rect 4512 4452 4540 4508
rect 4188 4428 4540 4452
rect 4188 4378 4216 4428
rect 4272 4378 4296 4428
rect 4352 4378 4376 4428
rect 4432 4378 4456 4428
rect 4512 4378 4540 4428
rect 4188 4326 4210 4378
rect 4272 4372 4274 4378
rect 4454 4372 4456 4378
rect 4262 4348 4274 4372
rect 4326 4348 4338 4372
rect 4390 4348 4402 4372
rect 4454 4348 4466 4372
rect 4272 4326 4274 4348
rect 4454 4326 4456 4348
rect 4518 4326 4540 4378
rect 4188 4292 4216 4326
rect 4272 4292 4296 4326
rect 4352 4292 4376 4326
rect 4432 4292 4456 4326
rect 4512 4292 4540 4326
rect 4188 3290 4540 4292
rect 4188 3238 4210 3290
rect 4262 3238 4274 3290
rect 4326 3238 4338 3290
rect 4390 3238 4402 3290
rect 4454 3238 4466 3290
rect 4518 3238 4540 3290
rect 4188 2202 4540 3238
rect 4188 2150 4210 2202
rect 4262 2150 4274 2202
rect 4326 2150 4338 2202
rect 4390 2150 4402 2202
rect 4454 2150 4466 2202
rect 4518 2150 4540 2202
rect 4188 1114 4540 2150
rect 4188 1062 4210 1114
rect 4262 1062 4274 1114
rect 4326 1062 4338 1114
rect 4390 1062 4402 1114
rect 4454 1062 4466 1114
rect 4518 1062 4540 1114
rect 4188 1040 4540 1062
rect 11836 4922 12188 5972
rect 11836 4870 11858 4922
rect 11910 4870 11922 4922
rect 11974 4870 11986 4922
rect 12038 4870 12050 4922
rect 12102 4870 12114 4922
rect 12166 4870 12188 4922
rect 11836 3834 12188 4870
rect 11836 3782 11858 3834
rect 11910 3782 11922 3834
rect 11974 3782 11986 3834
rect 12038 3782 12050 3834
rect 12102 3782 12114 3834
rect 12166 3782 12188 3834
rect 11836 2746 12188 3782
rect 11836 2694 11858 2746
rect 11910 2694 11922 2746
rect 11974 2694 11986 2746
rect 12038 2694 12050 2746
rect 12102 2694 12114 2746
rect 12166 2694 12188 2746
rect 11836 2236 12188 2694
rect 11836 2180 11864 2236
rect 11920 2180 11944 2236
rect 12000 2180 12024 2236
rect 12080 2180 12104 2236
rect 12160 2180 12188 2236
rect 11836 2156 12188 2180
rect 11836 2100 11864 2156
rect 11920 2100 11944 2156
rect 12000 2100 12024 2156
rect 12080 2100 12104 2156
rect 12160 2100 12188 2156
rect 11836 2076 12188 2100
rect 11836 2020 11864 2076
rect 11920 2020 11944 2076
rect 12000 2020 12024 2076
rect 12080 2020 12104 2076
rect 12160 2020 12188 2076
rect 11836 1996 12188 2020
rect 11836 1940 11864 1996
rect 11920 1940 11944 1996
rect 12000 1940 12024 1996
rect 12080 1940 12104 1996
rect 12160 1940 12188 1996
rect 11836 1658 12188 1940
rect 11836 1606 11858 1658
rect 11910 1606 11922 1658
rect 11974 1606 11986 1658
rect 12038 1606 12050 1658
rect 12102 1606 12114 1658
rect 12166 1606 12188 1658
rect 11836 1040 12188 1606
rect 14188 5466 14540 5972
rect 14188 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 14540 5466
rect 14188 4588 14540 5414
rect 14188 4532 14216 4588
rect 14272 4532 14296 4588
rect 14352 4532 14376 4588
rect 14432 4532 14456 4588
rect 14512 4532 14540 4588
rect 14188 4508 14540 4532
rect 14188 4452 14216 4508
rect 14272 4452 14296 4508
rect 14352 4452 14376 4508
rect 14432 4452 14456 4508
rect 14512 4452 14540 4508
rect 14188 4428 14540 4452
rect 14188 4378 14216 4428
rect 14272 4378 14296 4428
rect 14352 4378 14376 4428
rect 14432 4378 14456 4428
rect 14512 4378 14540 4428
rect 14188 4326 14210 4378
rect 14272 4372 14274 4378
rect 14454 4372 14456 4378
rect 14262 4348 14274 4372
rect 14326 4348 14338 4372
rect 14390 4348 14402 4372
rect 14454 4348 14466 4372
rect 14272 4326 14274 4348
rect 14454 4326 14456 4348
rect 14518 4326 14540 4378
rect 14188 4292 14216 4326
rect 14272 4292 14296 4326
rect 14352 4292 14376 4326
rect 14432 4292 14456 4326
rect 14512 4292 14540 4326
rect 14188 3290 14540 4292
rect 14188 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 14540 3290
rect 14188 2202 14540 3238
rect 14188 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 14540 2202
rect 14188 1114 14540 2150
rect 14188 1062 14210 1114
rect 14262 1062 14274 1114
rect 14326 1062 14338 1114
rect 14390 1062 14402 1114
rect 14454 1062 14466 1114
rect 14518 1062 14540 1114
rect 14188 1040 14540 1062
rect 21836 4922 22188 5972
rect 21836 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 21986 4922
rect 22038 4870 22050 4922
rect 22102 4870 22114 4922
rect 22166 4870 22188 4922
rect 21836 3834 22188 4870
rect 21836 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 21986 3834
rect 22038 3782 22050 3834
rect 22102 3782 22114 3834
rect 22166 3782 22188 3834
rect 21836 2746 22188 3782
rect 21836 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 21986 2746
rect 22038 2694 22050 2746
rect 22102 2694 22114 2746
rect 22166 2694 22188 2746
rect 21836 2236 22188 2694
rect 21836 2180 21864 2236
rect 21920 2180 21944 2236
rect 22000 2180 22024 2236
rect 22080 2180 22104 2236
rect 22160 2180 22188 2236
rect 21836 2156 22188 2180
rect 21836 2100 21864 2156
rect 21920 2100 21944 2156
rect 22000 2100 22024 2156
rect 22080 2100 22104 2156
rect 22160 2100 22188 2156
rect 21836 2076 22188 2100
rect 21836 2020 21864 2076
rect 21920 2020 21944 2076
rect 22000 2020 22024 2076
rect 22080 2020 22104 2076
rect 22160 2020 22188 2076
rect 21836 1996 22188 2020
rect 21836 1940 21864 1996
rect 21920 1940 21944 1996
rect 22000 1940 22024 1996
rect 22080 1940 22104 1996
rect 22160 1940 22188 1996
rect 21836 1658 22188 1940
rect 21836 1606 21858 1658
rect 21910 1606 21922 1658
rect 21974 1606 21986 1658
rect 22038 1606 22050 1658
rect 22102 1606 22114 1658
rect 22166 1606 22188 1658
rect 21836 1040 22188 1606
rect 24188 5466 24540 5972
rect 29828 5568 29880 5574
rect 29828 5510 29880 5516
rect 24188 5414 24210 5466
rect 24262 5414 24274 5466
rect 24326 5414 24338 5466
rect 24390 5414 24402 5466
rect 24454 5414 24466 5466
rect 24518 5414 24540 5466
rect 24188 4588 24540 5414
rect 24188 4532 24216 4588
rect 24272 4532 24296 4588
rect 24352 4532 24376 4588
rect 24432 4532 24456 4588
rect 24512 4532 24540 4588
rect 29368 4616 29420 4622
rect 29368 4558 29420 4564
rect 24188 4508 24540 4532
rect 24188 4452 24216 4508
rect 24272 4452 24296 4508
rect 24352 4452 24376 4508
rect 24432 4452 24456 4508
rect 24512 4452 24540 4508
rect 24188 4428 24540 4452
rect 24188 4378 24216 4428
rect 24272 4378 24296 4428
rect 24352 4378 24376 4428
rect 24432 4378 24456 4428
rect 24512 4378 24540 4428
rect 24188 4326 24210 4378
rect 24272 4372 24274 4378
rect 24454 4372 24456 4378
rect 24262 4348 24274 4372
rect 24326 4348 24338 4372
rect 24390 4348 24402 4372
rect 24454 4348 24466 4372
rect 24272 4326 24274 4348
rect 24454 4326 24456 4348
rect 24518 4326 24540 4378
rect 24188 4292 24216 4326
rect 24272 4292 24296 4326
rect 24352 4292 24376 4326
rect 24432 4292 24456 4326
rect 24512 4292 24540 4326
rect 24188 3290 24540 4292
rect 29380 4214 29408 4558
rect 29460 4548 29512 4554
rect 29460 4490 29512 4496
rect 29368 4208 29420 4214
rect 29368 4150 29420 4156
rect 28080 4072 28132 4078
rect 28080 4014 28132 4020
rect 29000 4072 29052 4078
rect 29000 4014 29052 4020
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 26896 3505 26924 3538
rect 27160 3528 27212 3534
rect 26882 3496 26938 3505
rect 26608 3460 26660 3466
rect 27160 3470 27212 3476
rect 26882 3431 26938 3440
rect 26608 3402 26660 3408
rect 24188 3238 24210 3290
rect 24262 3238 24274 3290
rect 24326 3238 24338 3290
rect 24390 3238 24402 3290
rect 24454 3238 24466 3290
rect 24518 3238 24540 3290
rect 24188 2202 24540 3238
rect 25688 3052 25740 3058
rect 25688 2994 25740 3000
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24188 2150 24210 2202
rect 24262 2150 24274 2202
rect 24326 2150 24338 2202
rect 24390 2150 24402 2202
rect 24454 2150 24466 2202
rect 24518 2150 24540 2202
rect 23940 1420 23992 1426
rect 23940 1362 23992 1368
rect 23480 1352 23532 1358
rect 23480 1294 23532 1300
rect 23032 870 23152 898
rect 23032 800 23060 870
rect 23018 0 23074 800
rect 23124 134 23152 870
rect 23492 800 23520 1294
rect 23952 800 23980 1362
rect 24188 1114 24540 2150
rect 24676 1964 24728 1970
rect 24676 1906 24728 1912
rect 24188 1062 24210 1114
rect 24262 1062 24274 1114
rect 24326 1062 24338 1114
rect 24390 1062 24402 1114
rect 24454 1062 24466 1114
rect 24518 1062 24540 1114
rect 24188 1040 24540 1062
rect 24412 870 24532 898
rect 24412 800 24440 870
rect 23112 128 23164 134
rect 23112 70 23164 76
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24398 0 24454 800
rect 24504 762 24532 870
rect 24688 762 24716 1906
rect 24872 800 24900 2382
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 25148 1494 25176 2246
rect 25240 1902 25268 2246
rect 25700 2106 25728 2994
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 25688 2100 25740 2106
rect 25688 2042 25740 2048
rect 25320 1964 25372 1970
rect 25320 1906 25372 1912
rect 25228 1896 25280 1902
rect 25228 1838 25280 1844
rect 25136 1488 25188 1494
rect 25136 1430 25188 1436
rect 25332 800 25360 1906
rect 25412 1896 25464 1902
rect 25412 1838 25464 1844
rect 25424 1562 25452 1838
rect 25412 1556 25464 1562
rect 25412 1498 25464 1504
rect 25688 1352 25740 1358
rect 25688 1294 25740 1300
rect 25700 1018 25728 1294
rect 25688 1012 25740 1018
rect 25688 954 25740 960
rect 26252 800 26280 2450
rect 26620 2106 26648 3402
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 26712 2106 26740 2994
rect 26884 2984 26936 2990
rect 26884 2926 26936 2932
rect 26792 2372 26844 2378
rect 26792 2314 26844 2320
rect 26608 2100 26660 2106
rect 26608 2042 26660 2048
rect 26700 2100 26752 2106
rect 26700 2042 26752 2048
rect 26804 1170 26832 2314
rect 26896 1358 26924 2926
rect 27172 2650 27200 3470
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 27068 2508 27120 2514
rect 27068 2450 27120 2456
rect 27080 2106 27108 2450
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 27068 2100 27120 2106
rect 27068 2042 27120 2048
rect 26884 1352 26936 1358
rect 26884 1294 26936 1300
rect 26712 1142 26832 1170
rect 26712 800 26740 1142
rect 27172 800 27200 2382
rect 27540 1902 27568 3878
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 27804 3392 27856 3398
rect 27804 3334 27856 3340
rect 27620 2372 27672 2378
rect 27620 2314 27672 2320
rect 27528 1896 27580 1902
rect 27528 1838 27580 1844
rect 27252 1352 27304 1358
rect 27252 1294 27304 1300
rect 27264 882 27292 1294
rect 27632 1222 27660 2314
rect 27816 1970 27844 3334
rect 28000 3194 28028 3470
rect 27988 3188 28040 3194
rect 27988 3130 28040 3136
rect 27804 1964 27856 1970
rect 27804 1906 27856 1912
rect 27620 1216 27672 1222
rect 27620 1158 27672 1164
rect 27252 876 27304 882
rect 27252 818 27304 824
rect 28092 800 28120 4014
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28644 3058 28672 3878
rect 28632 3052 28684 3058
rect 28632 2994 28684 3000
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 28184 1766 28212 2382
rect 28448 2304 28500 2310
rect 28448 2246 28500 2252
rect 28460 2106 28488 2246
rect 28448 2100 28500 2106
rect 28448 2042 28500 2048
rect 28172 1760 28224 1766
rect 28172 1702 28224 1708
rect 28264 1284 28316 1290
rect 28264 1226 28316 1232
rect 28540 1284 28592 1290
rect 28540 1226 28592 1232
rect 28276 1018 28304 1226
rect 28264 1012 28316 1018
rect 28264 954 28316 960
rect 28552 800 28580 1226
rect 29012 800 29040 4014
rect 29472 3194 29500 4490
rect 29840 4486 29868 5510
rect 29920 5092 29972 5098
rect 29920 5034 29972 5040
rect 29932 4690 29960 5034
rect 29920 4684 29972 4690
rect 29920 4626 29972 4632
rect 29828 4480 29880 4486
rect 29828 4422 29880 4428
rect 29932 4214 29960 4626
rect 29920 4208 29972 4214
rect 29920 4150 29972 4156
rect 29828 4072 29880 4078
rect 29826 4040 29828 4049
rect 29880 4040 29882 4049
rect 29826 3975 29882 3984
rect 29932 3602 29960 4150
rect 29920 3596 29972 3602
rect 29920 3538 29972 3544
rect 30300 3466 30328 6394
rect 30484 4554 30512 6462
rect 31024 6384 31076 6390
rect 31024 6326 31076 6332
rect 30746 5400 30802 5409
rect 31036 5370 31064 6326
rect 31574 6216 31630 6225
rect 31574 6151 31630 6160
rect 31116 5704 31168 5710
rect 31116 5646 31168 5652
rect 30746 5335 30802 5344
rect 31024 5364 31076 5370
rect 30760 5302 30788 5335
rect 31024 5306 31076 5312
rect 30748 5296 30800 5302
rect 30748 5238 30800 5244
rect 30564 5228 30616 5234
rect 30564 5170 30616 5176
rect 30472 4548 30524 4554
rect 30472 4490 30524 4496
rect 30484 4214 30512 4490
rect 30472 4208 30524 4214
rect 30472 4150 30524 4156
rect 30576 4026 30604 5170
rect 30760 4554 30788 5238
rect 30932 5228 30984 5234
rect 30932 5170 30984 5176
rect 30944 5137 30972 5170
rect 30930 5128 30986 5137
rect 30930 5063 30986 5072
rect 30840 5024 30892 5030
rect 30840 4966 30892 4972
rect 30748 4548 30800 4554
rect 30748 4490 30800 4496
rect 30656 4480 30708 4486
rect 30656 4422 30708 4428
rect 30668 4282 30696 4422
rect 30656 4276 30708 4282
rect 30656 4218 30708 4224
rect 30484 3998 30604 4026
rect 30656 4072 30708 4078
rect 30656 4014 30708 4020
rect 29736 3460 29788 3466
rect 29736 3402 29788 3408
rect 30288 3460 30340 3466
rect 30288 3402 30340 3408
rect 29460 3188 29512 3194
rect 29460 3130 29512 3136
rect 29092 2848 29144 2854
rect 29748 2825 29776 3402
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 29092 2790 29144 2796
rect 29734 2816 29790 2825
rect 29104 1970 29132 2790
rect 29734 2751 29790 2760
rect 29092 1964 29144 1970
rect 29092 1906 29144 1912
rect 29460 1556 29512 1562
rect 29460 1498 29512 1504
rect 29472 800 29500 1498
rect 29828 1352 29880 1358
rect 29828 1294 29880 1300
rect 29840 950 29868 1294
rect 29828 944 29880 950
rect 29828 886 29880 892
rect 29932 800 29960 2994
rect 30104 2984 30156 2990
rect 30104 2926 30156 2932
rect 30012 2916 30064 2922
rect 30012 2858 30064 2864
rect 30024 1358 30052 2858
rect 30116 2650 30144 2926
rect 30104 2644 30156 2650
rect 30104 2586 30156 2592
rect 30380 1896 30432 1902
rect 30380 1838 30432 1844
rect 30012 1352 30064 1358
rect 30012 1294 30064 1300
rect 30392 800 30420 1838
rect 30484 1494 30512 3998
rect 30668 3602 30696 4014
rect 30656 3596 30708 3602
rect 30656 3538 30708 3544
rect 30852 3058 30880 4966
rect 31036 4706 31064 5306
rect 31128 5302 31156 5646
rect 31392 5364 31444 5370
rect 31392 5306 31444 5312
rect 31116 5296 31168 5302
rect 31116 5238 31168 5244
rect 31208 5296 31260 5302
rect 31208 5238 31260 5244
rect 31220 4826 31248 5238
rect 31300 5228 31352 5234
rect 31300 5170 31352 5176
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 31312 4706 31340 5170
rect 31404 5030 31432 5306
rect 31392 5024 31444 5030
rect 31392 4966 31444 4972
rect 31036 4678 31156 4706
rect 30932 4616 30984 4622
rect 30932 4558 30984 4564
rect 30944 4146 30972 4558
rect 31128 4554 31156 4678
rect 31220 4678 31340 4706
rect 31116 4548 31168 4554
rect 31116 4490 31168 4496
rect 31024 4480 31076 4486
rect 31024 4422 31076 4428
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 31036 4078 31064 4422
rect 31024 4072 31076 4078
rect 31024 4014 31076 4020
rect 31024 3936 31076 3942
rect 31024 3878 31076 3884
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 30932 3460 30984 3466
rect 30932 3402 30984 3408
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 30576 2514 30604 2790
rect 30564 2508 30616 2514
rect 30564 2450 30616 2456
rect 30840 2440 30892 2446
rect 30562 2408 30618 2417
rect 30840 2382 30892 2388
rect 30562 2343 30618 2352
rect 30576 1766 30604 2343
rect 30564 1760 30616 1766
rect 30564 1702 30616 1708
rect 30472 1488 30524 1494
rect 30472 1430 30524 1436
rect 30852 1426 30880 2382
rect 30840 1420 30892 1426
rect 30840 1362 30892 1368
rect 30840 1012 30892 1018
rect 30840 954 30892 960
rect 30852 800 30880 954
rect 24504 734 24716 762
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26238 0 26294 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 30944 746 30972 3402
rect 31036 3126 31064 3878
rect 31024 3120 31076 3126
rect 31024 3062 31076 3068
rect 31128 2972 31156 3878
rect 31036 2944 31156 2972
rect 31036 2854 31064 2944
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 31220 2774 31248 4678
rect 31588 4570 31616 6151
rect 31666 5264 31722 5273
rect 31666 5199 31668 5208
rect 31720 5199 31722 5208
rect 31668 5170 31720 5176
rect 31836 4922 32188 5972
rect 32416 5358 32628 5386
rect 32416 5302 32444 5358
rect 32600 5302 32628 5358
rect 32404 5296 32456 5302
rect 32218 5264 32274 5273
rect 32588 5296 32640 5302
rect 32404 5238 32456 5244
rect 32494 5264 32550 5273
rect 32218 5199 32274 5208
rect 32588 5238 32640 5244
rect 32494 5199 32496 5208
rect 32232 5098 32260 5199
rect 32548 5199 32550 5208
rect 32496 5170 32548 5176
rect 32312 5160 32364 5166
rect 32404 5160 32456 5166
rect 32312 5102 32364 5108
rect 32402 5128 32404 5137
rect 32456 5128 32458 5137
rect 32220 5092 32272 5098
rect 32220 5034 32272 5040
rect 31836 4870 31858 4922
rect 31910 4870 31922 4922
rect 31974 4870 31986 4922
rect 32038 4870 32050 4922
rect 32102 4870 32114 4922
rect 32166 4870 32188 4922
rect 31588 4542 31708 4570
rect 31300 4480 31352 4486
rect 31300 4422 31352 4428
rect 31312 4282 31340 4422
rect 31300 4276 31352 4282
rect 31352 4236 31432 4264
rect 31300 4218 31352 4224
rect 31404 3602 31432 4236
rect 31680 4078 31708 4542
rect 31668 4072 31720 4078
rect 31668 4014 31720 4020
rect 31680 3942 31708 4014
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 31836 3834 32188 4870
rect 32324 4758 32352 5102
rect 32402 5063 32458 5072
rect 32402 4992 32458 5001
rect 32402 4927 32458 4936
rect 32416 4826 32444 4927
rect 32404 4820 32456 4826
rect 32404 4762 32456 4768
rect 32312 4752 32364 4758
rect 32312 4694 32364 4700
rect 32324 4298 32352 4694
rect 32324 4270 32444 4298
rect 32310 4176 32366 4185
rect 32310 4111 32366 4120
rect 32324 4078 32352 4111
rect 32312 4072 32364 4078
rect 32312 4014 32364 4020
rect 32220 3936 32272 3942
rect 32220 3878 32272 3884
rect 31836 3782 31858 3834
rect 31910 3782 31922 3834
rect 31974 3782 31986 3834
rect 32038 3782 32050 3834
rect 32102 3782 32114 3834
rect 32166 3782 32188 3834
rect 31693 3664 31745 3670
rect 31680 3612 31693 3652
rect 31680 3606 31745 3612
rect 31392 3596 31444 3602
rect 31392 3538 31444 3544
rect 31484 3596 31536 3602
rect 31484 3538 31536 3544
rect 31404 3398 31432 3538
rect 31392 3392 31444 3398
rect 31392 3334 31444 3340
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31312 2854 31340 3130
rect 31496 3058 31524 3538
rect 31680 3233 31708 3606
rect 31666 3224 31722 3233
rect 31666 3159 31722 3168
rect 31484 3052 31536 3058
rect 31484 2994 31536 3000
rect 31668 2984 31720 2990
rect 31720 2944 31800 2972
rect 31668 2926 31720 2932
rect 31300 2848 31352 2854
rect 31300 2790 31352 2796
rect 31128 2746 31248 2774
rect 31128 1970 31156 2746
rect 31484 2440 31536 2446
rect 31484 2382 31536 2388
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31116 1964 31168 1970
rect 31116 1906 31168 1912
rect 31312 800 31340 2246
rect 31496 1562 31524 2382
rect 31484 1556 31536 1562
rect 31484 1498 31536 1504
rect 31772 800 31800 2944
rect 31836 2746 32188 3782
rect 32232 3097 32260 3878
rect 32324 3738 32352 4014
rect 32416 3942 32444 4270
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 32312 3732 32364 3738
rect 32312 3674 32364 3680
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 32416 3369 32444 3606
rect 32402 3360 32458 3369
rect 32402 3295 32458 3304
rect 32218 3088 32274 3097
rect 32218 3023 32274 3032
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 31836 2694 31858 2746
rect 31910 2694 31922 2746
rect 31974 2694 31986 2746
rect 32038 2694 32050 2746
rect 32102 2694 32114 2746
rect 32166 2694 32188 2746
rect 31836 2236 32188 2694
rect 32232 2650 32260 2926
rect 32220 2644 32272 2650
rect 32220 2586 32272 2592
rect 32508 2514 32536 5170
rect 32772 4616 32824 4622
rect 32772 4558 32824 4564
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 32588 4004 32640 4010
rect 32640 3964 32720 3992
rect 32588 3946 32640 3952
rect 32586 3632 32642 3641
rect 32586 3567 32642 3576
rect 32600 3534 32628 3567
rect 32588 3528 32640 3534
rect 32588 3470 32640 3476
rect 32600 3194 32628 3470
rect 32588 3188 32640 3194
rect 32588 3130 32640 3136
rect 32496 2508 32548 2514
rect 32496 2450 32548 2456
rect 32496 2304 32548 2310
rect 32496 2246 32548 2252
rect 31836 2180 31864 2236
rect 31920 2180 31944 2236
rect 32000 2180 32024 2236
rect 32080 2180 32104 2236
rect 32160 2180 32188 2236
rect 31836 2156 32188 2180
rect 31836 2100 31864 2156
rect 31920 2100 31944 2156
rect 32000 2100 32024 2156
rect 32080 2100 32104 2156
rect 32160 2100 32188 2156
rect 31836 2076 32188 2100
rect 31836 2020 31864 2076
rect 31920 2020 31944 2076
rect 32000 2020 32024 2076
rect 32080 2020 32104 2076
rect 32160 2020 32188 2076
rect 31836 1996 32188 2020
rect 31836 1940 31864 1996
rect 31920 1940 31944 1996
rect 32000 1940 32024 1996
rect 32080 1940 32104 1996
rect 32160 1940 32188 1996
rect 31836 1658 32188 1940
rect 32220 1896 32272 1902
rect 32220 1838 32272 1844
rect 31836 1606 31858 1658
rect 31910 1606 31922 1658
rect 31974 1606 31986 1658
rect 32038 1606 32050 1658
rect 32102 1606 32114 1658
rect 32166 1606 32188 1658
rect 31836 1040 32188 1606
rect 32232 800 32260 1838
rect 32508 1766 32536 2246
rect 32496 1760 32548 1766
rect 32496 1702 32548 1708
rect 32692 1494 32720 3964
rect 32784 3194 32812 4558
rect 32772 3188 32824 3194
rect 32772 3130 32824 3136
rect 32876 1562 32904 4558
rect 32968 4486 32996 7550
rect 35164 6724 35216 6730
rect 35164 6666 35216 6672
rect 33692 6588 33744 6594
rect 33692 6530 33744 6536
rect 33232 5636 33284 5642
rect 33232 5578 33284 5584
rect 32956 4480 33008 4486
rect 32956 4422 33008 4428
rect 32968 4214 32996 4422
rect 32956 4208 33008 4214
rect 32956 4150 33008 4156
rect 32956 4072 33008 4078
rect 32956 4014 33008 4020
rect 32968 3670 32996 4014
rect 33140 3936 33192 3942
rect 33140 3878 33192 3884
rect 32956 3664 33008 3670
rect 32956 3606 33008 3612
rect 32968 3466 32996 3606
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 32956 3460 33008 3466
rect 32956 3402 33008 3408
rect 33060 1970 33088 3538
rect 33152 2990 33180 3878
rect 33140 2984 33192 2990
rect 33140 2926 33192 2932
rect 33140 2848 33192 2854
rect 33244 2802 33272 5578
rect 33600 4480 33652 4486
rect 33600 4422 33652 4428
rect 33612 4282 33640 4422
rect 33600 4276 33652 4282
rect 33600 4218 33652 4224
rect 33598 4176 33654 4185
rect 33598 4111 33654 4120
rect 33324 4072 33376 4078
rect 33324 4014 33376 4020
rect 33336 3738 33364 4014
rect 33508 3936 33560 3942
rect 33414 3904 33470 3913
rect 33508 3878 33560 3884
rect 33414 3839 33470 3848
rect 33324 3732 33376 3738
rect 33324 3674 33376 3680
rect 33324 3528 33376 3534
rect 33428 3516 33456 3839
rect 33376 3488 33456 3516
rect 33324 3470 33376 3476
rect 33416 3392 33468 3398
rect 33416 3334 33468 3340
rect 33324 3120 33376 3126
rect 33324 3062 33376 3068
rect 33192 2796 33272 2802
rect 33140 2790 33272 2796
rect 33152 2774 33272 2790
rect 33048 1964 33100 1970
rect 33048 1906 33100 1912
rect 32864 1556 32916 1562
rect 32864 1498 32916 1504
rect 32680 1488 32732 1494
rect 32680 1430 32732 1436
rect 33140 1420 33192 1426
rect 33140 1362 33192 1368
rect 32600 882 32720 898
rect 32588 876 32720 882
rect 32640 870 32720 876
rect 32588 818 32640 824
rect 32692 800 32720 870
rect 33152 800 33180 1362
rect 33336 1018 33364 3062
rect 33428 2961 33456 3334
rect 33414 2952 33470 2961
rect 33414 2887 33470 2896
rect 33416 2848 33468 2854
rect 33416 2790 33468 2796
rect 33324 1012 33376 1018
rect 33324 954 33376 960
rect 33428 814 33456 2790
rect 33520 1970 33548 3878
rect 33612 3398 33640 4111
rect 33704 4078 33732 6530
rect 33782 6352 33838 6361
rect 33782 6287 33838 6296
rect 33692 4072 33744 4078
rect 33692 4014 33744 4020
rect 33796 3942 33824 6287
rect 34188 5466 34540 5972
rect 34796 5704 34848 5710
rect 34796 5646 34848 5652
rect 34188 5414 34210 5466
rect 34262 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 34540 5466
rect 34058 5128 34114 5137
rect 34058 5063 34114 5072
rect 33966 4856 34022 4865
rect 34072 4826 34100 5063
rect 33966 4791 34022 4800
rect 34060 4820 34112 4826
rect 33980 4690 34008 4791
rect 34060 4762 34112 4768
rect 33968 4684 34020 4690
rect 33968 4626 34020 4632
rect 34188 4588 34540 5414
rect 34612 5228 34664 5234
rect 34612 5170 34664 5176
rect 34624 4622 34652 5170
rect 34704 5024 34756 5030
rect 34704 4966 34756 4972
rect 34716 4865 34744 4966
rect 34702 4856 34758 4865
rect 34702 4791 34758 4800
rect 33876 4548 33928 4554
rect 33876 4490 33928 4496
rect 33968 4548 34020 4554
rect 33968 4490 34020 4496
rect 34188 4532 34216 4588
rect 34272 4532 34296 4588
rect 34352 4532 34376 4588
rect 34432 4532 34456 4588
rect 34512 4532 34540 4588
rect 34612 4616 34664 4622
rect 34808 4604 34836 5646
rect 34886 5400 34942 5409
rect 34886 5335 34942 5344
rect 34612 4558 34664 4564
rect 34716 4576 34836 4604
rect 34188 4508 34540 4532
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33796 3754 33824 3878
rect 33704 3726 33824 3754
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33704 3194 33732 3726
rect 33782 3360 33838 3369
rect 33782 3295 33838 3304
rect 33796 3194 33824 3295
rect 33692 3188 33744 3194
rect 33692 3130 33744 3136
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33888 2650 33916 4490
rect 33980 4214 34008 4490
rect 34188 4452 34216 4508
rect 34272 4452 34296 4508
rect 34352 4452 34376 4508
rect 34432 4452 34456 4508
rect 34512 4452 34540 4508
rect 34188 4428 34540 4452
rect 34188 4378 34216 4428
rect 34272 4378 34296 4428
rect 34352 4378 34376 4428
rect 34432 4378 34456 4428
rect 34512 4378 34540 4428
rect 34188 4326 34210 4378
rect 34272 4372 34274 4378
rect 34454 4372 34456 4378
rect 34262 4348 34274 4372
rect 34326 4348 34338 4372
rect 34390 4348 34402 4372
rect 34454 4348 34466 4372
rect 34272 4326 34274 4348
rect 34454 4326 34456 4348
rect 34518 4326 34540 4378
rect 34188 4292 34216 4326
rect 34272 4292 34296 4326
rect 34352 4292 34376 4326
rect 34432 4292 34456 4326
rect 34512 4292 34540 4326
rect 34060 4276 34112 4282
rect 34060 4218 34112 4224
rect 33968 4208 34020 4214
rect 34072 4185 34100 4218
rect 33968 4150 34020 4156
rect 34058 4176 34114 4185
rect 34058 4111 34114 4120
rect 34060 4072 34112 4078
rect 33980 4032 34060 4060
rect 33980 3777 34008 4032
rect 34060 4014 34112 4020
rect 34060 3936 34112 3942
rect 34060 3878 34112 3884
rect 33966 3768 34022 3777
rect 33966 3703 34022 3712
rect 33980 3670 34008 3703
rect 33968 3664 34020 3670
rect 33968 3606 34020 3612
rect 33980 3534 34008 3606
rect 33968 3528 34020 3534
rect 33968 3470 34020 3476
rect 34072 3466 34100 3878
rect 34060 3460 34112 3466
rect 34060 3402 34112 3408
rect 33968 3392 34020 3398
rect 33966 3360 33968 3369
rect 34020 3360 34022 3369
rect 33966 3295 34022 3304
rect 34188 3290 34540 4292
rect 34716 4214 34744 4576
rect 34900 4282 34928 5335
rect 35176 5030 35204 6666
rect 35900 5704 35952 5710
rect 35900 5646 35952 5652
rect 35806 5400 35862 5409
rect 35806 5335 35862 5344
rect 35622 5128 35678 5137
rect 35622 5063 35678 5072
rect 35164 5024 35216 5030
rect 35164 4966 35216 4972
rect 35532 5024 35584 5030
rect 35532 4966 35584 4972
rect 34978 4856 35034 4865
rect 34978 4791 35034 4800
rect 34992 4690 35020 4791
rect 34980 4684 35032 4690
rect 34980 4626 35032 4632
rect 35164 4616 35216 4622
rect 35216 4576 35296 4604
rect 35164 4558 35216 4564
rect 35072 4548 35124 4554
rect 35072 4490 35124 4496
rect 34888 4276 34940 4282
rect 34888 4218 34940 4224
rect 34980 4276 35032 4282
rect 34980 4218 35032 4224
rect 34704 4208 34756 4214
rect 34704 4150 34756 4156
rect 34992 4128 35020 4218
rect 34900 4100 35020 4128
rect 34796 4072 34848 4078
rect 34796 4014 34848 4020
rect 34808 3738 34836 4014
rect 34796 3732 34848 3738
rect 34796 3674 34848 3680
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34188 3238 34210 3290
rect 34262 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 34540 3290
rect 34060 3120 34112 3126
rect 34060 3062 34112 3068
rect 33876 2644 33928 2650
rect 33876 2586 33928 2592
rect 33874 2544 33930 2553
rect 33600 2508 33652 2514
rect 33874 2479 33930 2488
rect 33600 2450 33652 2456
rect 33508 1964 33560 1970
rect 33508 1906 33560 1912
rect 33416 808 33468 814
rect 30932 740 30984 746
rect 30932 682 30984 688
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32678 0 32734 800
rect 33138 0 33194 800
rect 33612 800 33640 2450
rect 33888 1970 33916 2479
rect 33968 2440 34020 2446
rect 33968 2382 34020 2388
rect 33980 2038 34008 2382
rect 34072 2106 34100 3062
rect 34188 2202 34540 3238
rect 34188 2150 34210 2202
rect 34262 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 34540 2202
rect 34060 2100 34112 2106
rect 34060 2042 34112 2048
rect 33968 2032 34020 2038
rect 33968 1974 34020 1980
rect 33876 1964 33928 1970
rect 33876 1906 33928 1912
rect 34060 1896 34112 1902
rect 34060 1838 34112 1844
rect 33968 1352 34020 1358
rect 33966 1320 33968 1329
rect 34020 1320 34022 1329
rect 33966 1255 34022 1264
rect 34072 800 34100 1838
rect 34188 1114 34540 2150
rect 34624 1970 34652 3334
rect 34900 2417 34928 4100
rect 35084 3890 35112 4490
rect 35164 4480 35216 4486
rect 35164 4422 35216 4428
rect 35176 4185 35204 4422
rect 35268 4264 35296 4576
rect 35348 4276 35400 4282
rect 35268 4236 35348 4264
rect 35348 4218 35400 4224
rect 35440 4208 35492 4214
rect 35162 4176 35218 4185
rect 35162 4111 35218 4120
rect 35438 4176 35440 4185
rect 35492 4176 35494 4185
rect 35544 4146 35572 4966
rect 35636 4486 35664 5063
rect 35716 4616 35768 4622
rect 35716 4558 35768 4564
rect 35624 4480 35676 4486
rect 35624 4422 35676 4428
rect 35728 4146 35756 4558
rect 35820 4282 35848 5335
rect 35808 4276 35860 4282
rect 35808 4218 35860 4224
rect 35912 4214 35940 5646
rect 35900 4208 35952 4214
rect 35900 4150 35952 4156
rect 35438 4111 35494 4120
rect 35532 4140 35584 4146
rect 35176 4026 35204 4111
rect 35532 4082 35584 4088
rect 35716 4140 35768 4146
rect 35716 4082 35768 4088
rect 35808 4140 35860 4146
rect 35808 4082 35860 4088
rect 35176 3998 35388 4026
rect 35544 4010 35572 4082
rect 35084 3862 35204 3890
rect 34980 3392 35032 3398
rect 34978 3360 34980 3369
rect 35072 3392 35124 3398
rect 35032 3360 35034 3369
rect 35072 3334 35124 3340
rect 34978 3295 35034 3304
rect 35084 2922 35112 3334
rect 35072 2916 35124 2922
rect 35072 2858 35124 2864
rect 34980 2440 35032 2446
rect 34886 2408 34942 2417
rect 34980 2382 35032 2388
rect 34886 2343 34942 2352
rect 34888 2032 34940 2038
rect 34888 1974 34940 1980
rect 34612 1964 34664 1970
rect 34612 1906 34664 1912
rect 34900 1494 34928 1974
rect 34888 1488 34940 1494
rect 34888 1430 34940 1436
rect 34188 1062 34210 1114
rect 34262 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 34540 1114
rect 34188 1040 34540 1062
rect 34520 944 34572 950
rect 34520 886 34572 892
rect 34532 800 34560 886
rect 34992 800 35020 2382
rect 35176 2310 35204 3862
rect 35254 3768 35310 3777
rect 35254 3703 35310 3712
rect 35268 3602 35296 3703
rect 35256 3596 35308 3602
rect 35256 3538 35308 3544
rect 35360 3466 35388 3998
rect 35440 4004 35492 4010
rect 35440 3946 35492 3952
rect 35532 4004 35584 4010
rect 35532 3946 35584 3952
rect 35452 3466 35480 3946
rect 35348 3460 35400 3466
rect 35348 3402 35400 3408
rect 35440 3460 35492 3466
rect 35440 3402 35492 3408
rect 35544 3398 35572 3946
rect 35728 3777 35756 4082
rect 35714 3768 35770 3777
rect 35714 3703 35770 3712
rect 35532 3392 35584 3398
rect 35532 3334 35584 3340
rect 35716 3392 35768 3398
rect 35716 3334 35768 3340
rect 35532 3120 35584 3126
rect 35532 3062 35584 3068
rect 35544 2972 35572 3062
rect 35728 2972 35756 3334
rect 35438 2952 35494 2961
rect 35544 2944 35756 2972
rect 35438 2887 35494 2896
rect 35164 2304 35216 2310
rect 35164 2246 35216 2252
rect 35452 1358 35480 2887
rect 35624 1896 35676 1902
rect 35624 1838 35676 1844
rect 35636 1562 35664 1838
rect 35820 1766 35848 4082
rect 36004 3738 36032 7686
rect 36084 7676 36136 7682
rect 36084 7618 36136 7624
rect 35992 3732 36044 3738
rect 35992 3674 36044 3680
rect 36096 3670 36124 7618
rect 48136 6860 48188 6866
rect 48136 6802 48188 6808
rect 36636 6792 36688 6798
rect 36636 6734 36688 6740
rect 36176 5568 36228 5574
rect 36176 5510 36228 5516
rect 36188 4622 36216 5510
rect 36452 5364 36504 5370
rect 36452 5306 36504 5312
rect 36464 5030 36492 5306
rect 36452 5024 36504 5030
rect 36266 4992 36322 5001
rect 36452 4966 36504 4972
rect 36266 4927 36322 4936
rect 36280 4690 36308 4927
rect 36268 4684 36320 4690
rect 36268 4626 36320 4632
rect 36176 4616 36228 4622
rect 36176 4558 36228 4564
rect 36648 4146 36676 6734
rect 40222 6488 40278 6497
rect 40222 6423 40278 6432
rect 37922 5264 37978 5273
rect 37922 5199 37978 5208
rect 36636 4140 36688 4146
rect 36636 4082 36688 4088
rect 36268 4072 36320 4078
rect 36268 4014 36320 4020
rect 36176 3936 36228 3942
rect 36280 3913 36308 4014
rect 36452 4004 36504 4010
rect 36452 3946 36504 3952
rect 36176 3878 36228 3884
rect 36266 3904 36322 3913
rect 36084 3664 36136 3670
rect 36084 3606 36136 3612
rect 36082 3224 36138 3233
rect 36082 3159 36138 3168
rect 35900 2984 35952 2990
rect 35900 2926 35952 2932
rect 35808 1760 35860 1766
rect 35808 1702 35860 1708
rect 35624 1556 35676 1562
rect 35624 1498 35676 1504
rect 35440 1352 35492 1358
rect 35440 1294 35492 1300
rect 35624 1284 35676 1290
rect 35624 1226 35676 1232
rect 35636 898 35664 1226
rect 35452 870 35664 898
rect 35452 800 35480 870
rect 35912 800 35940 2926
rect 36096 2854 36124 3159
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36084 2848 36136 2854
rect 36188 2825 36216 3878
rect 36266 3839 36322 3848
rect 36360 3528 36412 3534
rect 36360 3470 36412 3476
rect 36084 2790 36136 2796
rect 36174 2816 36230 2825
rect 36004 2514 36032 2790
rect 36174 2751 36230 2760
rect 36372 2650 36400 3470
rect 36464 3097 36492 3946
rect 36648 3777 36676 4082
rect 36634 3768 36690 3777
rect 36634 3703 36690 3712
rect 36544 3460 36596 3466
rect 36544 3402 36596 3408
rect 36450 3088 36506 3097
rect 36450 3023 36506 3032
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 35992 2508 36044 2514
rect 35992 2450 36044 2456
rect 36556 2106 36584 3402
rect 37462 3088 37518 3097
rect 37462 3023 37518 3032
rect 37648 3052 37700 3058
rect 37476 2990 37504 3023
rect 37648 2994 37700 3000
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 37660 2650 37688 2994
rect 37936 2990 37964 5199
rect 40040 4684 40092 4690
rect 40040 4626 40092 4632
rect 38384 3460 38436 3466
rect 38384 3402 38436 3408
rect 38396 3058 38424 3402
rect 38844 3392 38896 3398
rect 38844 3334 38896 3340
rect 38856 3058 38884 3334
rect 39764 3188 39816 3194
rect 39764 3130 39816 3136
rect 38200 3052 38252 3058
rect 38200 2994 38252 3000
rect 38384 3052 38436 3058
rect 38384 2994 38436 3000
rect 38844 3052 38896 3058
rect 38844 2994 38896 3000
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 37832 2984 37884 2990
rect 37832 2926 37884 2932
rect 37924 2984 37976 2990
rect 37924 2926 37976 2932
rect 37844 2650 37872 2926
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 37004 2440 37056 2446
rect 37004 2382 37056 2388
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 37016 2106 37044 2382
rect 36544 2100 36596 2106
rect 36544 2042 36596 2048
rect 37004 2100 37056 2106
rect 37004 2042 37056 2048
rect 37280 1896 37332 1902
rect 37280 1838 37332 1844
rect 36820 1828 36872 1834
rect 36820 1770 36872 1776
rect 36360 1352 36412 1358
rect 36360 1294 36412 1300
rect 36372 800 36400 1294
rect 36832 800 36860 1770
rect 37292 800 37320 1838
rect 37752 800 37780 2382
rect 38212 1358 38240 2994
rect 39132 2650 39160 2994
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 38752 2440 38804 2446
rect 38752 2382 38804 2388
rect 38764 1562 38792 2382
rect 39120 1896 39172 1902
rect 39120 1838 39172 1844
rect 38752 1556 38804 1562
rect 38752 1498 38804 1504
rect 38200 1352 38252 1358
rect 38200 1294 38252 1300
rect 38660 1352 38712 1358
rect 38660 1294 38712 1300
rect 38292 1284 38344 1290
rect 38292 1226 38344 1232
rect 38304 898 38332 1226
rect 38212 870 38332 898
rect 38212 800 38240 870
rect 38672 800 38700 1294
rect 39132 800 39160 1838
rect 39776 1358 39804 3130
rect 40052 1902 40080 4626
rect 40236 4078 40264 6423
rect 47308 6180 47360 6186
rect 47308 6122 47360 6128
rect 41512 5704 41564 5710
rect 41512 5646 41564 5652
rect 40776 4276 40828 4282
rect 40776 4218 40828 4224
rect 40788 4078 40816 4218
rect 40868 4140 40920 4146
rect 40868 4082 40920 4088
rect 40224 4072 40276 4078
rect 40224 4014 40276 4020
rect 40776 4072 40828 4078
rect 40776 4014 40828 4020
rect 40132 3596 40184 3602
rect 40132 3538 40184 3544
rect 40144 3346 40172 3538
rect 40236 3466 40264 4014
rect 40880 3738 40908 4082
rect 40960 4004 41012 4010
rect 40960 3946 41012 3952
rect 40868 3732 40920 3738
rect 40868 3674 40920 3680
rect 40224 3460 40276 3466
rect 40224 3402 40276 3408
rect 40316 3460 40368 3466
rect 40316 3402 40368 3408
rect 40328 3346 40356 3402
rect 40144 3318 40356 3346
rect 40972 2990 41000 3946
rect 41328 3732 41380 3738
rect 41328 3674 41380 3680
rect 41340 3058 41368 3674
rect 41524 3466 41552 5646
rect 41836 4922 42188 5972
rect 42708 5840 42760 5846
rect 42708 5782 42760 5788
rect 42524 5704 42576 5710
rect 42720 5681 42748 5782
rect 42524 5646 42576 5652
rect 42706 5672 42762 5681
rect 41836 4870 41858 4922
rect 41910 4870 41922 4922
rect 41974 4870 41986 4922
rect 42038 4870 42050 4922
rect 42102 4870 42114 4922
rect 42166 4870 42188 4922
rect 41836 3834 42188 4870
rect 42536 4078 42564 5646
rect 42706 5607 42762 5616
rect 44188 5466 44540 5972
rect 44732 5840 44784 5846
rect 44730 5808 44732 5817
rect 44784 5808 44786 5817
rect 44730 5743 44786 5752
rect 45560 5704 45612 5710
rect 45560 5646 45612 5652
rect 44188 5414 44210 5466
rect 44262 5414 44274 5466
rect 44326 5414 44338 5466
rect 44390 5414 44402 5466
rect 44454 5414 44466 5466
rect 44518 5414 44540 5466
rect 43904 5160 43956 5166
rect 43904 5102 43956 5108
rect 43916 5030 43944 5102
rect 43904 5024 43956 5030
rect 43904 4966 43956 4972
rect 44188 4588 44540 5414
rect 45284 5364 45336 5370
rect 45284 5306 45336 5312
rect 45376 5364 45428 5370
rect 45376 5306 45428 5312
rect 44916 5160 44968 5166
rect 44916 5102 44968 5108
rect 44188 4532 44216 4588
rect 44272 4532 44296 4588
rect 44352 4532 44376 4588
rect 44432 4532 44456 4588
rect 44512 4532 44540 4588
rect 44732 4616 44784 4622
rect 44732 4558 44784 4564
rect 44188 4508 44540 4532
rect 44188 4452 44216 4508
rect 44272 4452 44296 4508
rect 44352 4452 44376 4508
rect 44432 4452 44456 4508
rect 44512 4452 44540 4508
rect 44188 4428 44540 4452
rect 44188 4378 44216 4428
rect 44272 4378 44296 4428
rect 44352 4378 44376 4428
rect 44432 4378 44456 4428
rect 44512 4378 44540 4428
rect 44188 4326 44210 4378
rect 44272 4372 44274 4378
rect 44454 4372 44456 4378
rect 44262 4348 44274 4372
rect 44326 4348 44338 4372
rect 44390 4348 44402 4372
rect 44454 4348 44466 4372
rect 44272 4326 44274 4348
rect 44454 4326 44456 4348
rect 44518 4326 44540 4378
rect 44188 4292 44216 4326
rect 44272 4292 44296 4326
rect 44352 4292 44376 4326
rect 44432 4292 44456 4326
rect 44512 4292 44540 4326
rect 42340 4072 42392 4078
rect 42340 4014 42392 4020
rect 42524 4072 42576 4078
rect 42524 4014 42576 4020
rect 41836 3782 41858 3834
rect 41910 3782 41922 3834
rect 41974 3782 41986 3834
rect 42038 3782 42050 3834
rect 42102 3782 42114 3834
rect 42166 3782 42188 3834
rect 41512 3460 41564 3466
rect 41512 3402 41564 3408
rect 41604 3460 41656 3466
rect 41604 3402 41656 3408
rect 41328 3052 41380 3058
rect 41328 2994 41380 3000
rect 40960 2984 41012 2990
rect 40960 2926 41012 2932
rect 41616 2650 41644 3402
rect 41696 3052 41748 3058
rect 41696 2994 41748 3000
rect 41708 2650 41736 2994
rect 41836 2746 42188 3782
rect 42248 3460 42300 3466
rect 42248 3402 42300 3408
rect 42260 3194 42288 3402
rect 42248 3188 42300 3194
rect 42248 3130 42300 3136
rect 42248 2984 42300 2990
rect 42248 2926 42300 2932
rect 41836 2694 41858 2746
rect 41910 2694 41922 2746
rect 41974 2694 41986 2746
rect 42038 2694 42050 2746
rect 42102 2694 42114 2746
rect 42166 2694 42188 2746
rect 41604 2644 41656 2650
rect 41604 2586 41656 2592
rect 41696 2644 41748 2650
rect 41696 2586 41748 2592
rect 40684 2440 40736 2446
rect 40684 2382 40736 2388
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 40696 2106 40724 2382
rect 41432 2106 41460 2382
rect 41836 2236 42188 2694
rect 41836 2180 41864 2236
rect 41920 2180 41944 2236
rect 42000 2180 42024 2236
rect 42080 2180 42104 2236
rect 42160 2180 42188 2236
rect 41836 2156 42188 2180
rect 40684 2100 40736 2106
rect 40684 2042 40736 2048
rect 41420 2100 41472 2106
rect 41420 2042 41472 2048
rect 41696 2100 41748 2106
rect 41696 2042 41748 2048
rect 41836 2100 41864 2156
rect 41920 2100 41944 2156
rect 42000 2100 42024 2156
rect 42080 2100 42104 2156
rect 42160 2100 42188 2156
rect 41836 2076 42188 2100
rect 41144 2032 41196 2038
rect 41144 1974 41196 1980
rect 40040 1896 40092 1902
rect 40040 1838 40092 1844
rect 41156 1737 41184 1974
rect 41236 1964 41288 1970
rect 41236 1906 41288 1912
rect 41420 1964 41472 1970
rect 41420 1906 41472 1912
rect 41142 1728 41198 1737
rect 41142 1663 41198 1672
rect 41248 1562 41276 1906
rect 41236 1556 41288 1562
rect 41236 1498 41288 1504
rect 41432 1426 41460 1906
rect 41708 1766 41736 2042
rect 41836 2020 41864 2076
rect 41920 2020 41944 2076
rect 42000 2020 42024 2076
rect 42080 2020 42104 2076
rect 42160 2020 42188 2076
rect 41836 1996 42188 2020
rect 41836 1940 41864 1996
rect 41920 1940 41944 1996
rect 42000 1940 42024 1996
rect 42080 1940 42104 1996
rect 42160 1940 42188 1996
rect 41696 1760 41748 1766
rect 41696 1702 41748 1708
rect 41836 1658 42188 1940
rect 41836 1606 41858 1658
rect 41910 1606 41922 1658
rect 41974 1606 41986 1658
rect 42038 1606 42050 1658
rect 42102 1606 42114 1658
rect 42166 1606 42188 1658
rect 40500 1420 40552 1426
rect 40500 1362 40552 1368
rect 41420 1420 41472 1426
rect 41420 1362 41472 1368
rect 39764 1352 39816 1358
rect 39764 1294 39816 1300
rect 40040 1352 40092 1358
rect 40040 1294 40092 1300
rect 39580 1284 39632 1290
rect 39580 1226 39632 1232
rect 39592 800 39620 1226
rect 40052 800 40080 1294
rect 40512 800 40540 1362
rect 40960 1284 41012 1290
rect 40960 1226 41012 1232
rect 40972 800 41000 1226
rect 41836 1040 42188 1606
rect 41420 1012 41472 1018
rect 41420 954 41472 960
rect 41432 800 41460 954
rect 41892 870 42012 898
rect 41892 800 41920 870
rect 33416 750 33468 756
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34518 0 34574 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39118 0 39174 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 40958 0 41014 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 41984 762 42012 870
rect 42260 762 42288 2926
rect 42352 1358 42380 4014
rect 44188 3290 44540 4292
rect 44188 3238 44210 3290
rect 44262 3238 44274 3290
rect 44326 3238 44338 3290
rect 44390 3238 44402 3290
rect 44454 3238 44466 3290
rect 44518 3238 44540 3290
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 42444 2650 42472 2994
rect 42524 2848 42576 2854
rect 42524 2790 42576 2796
rect 42984 2848 43036 2854
rect 42984 2790 43036 2796
rect 42432 2644 42484 2650
rect 42432 2586 42484 2592
rect 42536 1970 42564 2790
rect 42996 2514 43024 2790
rect 42984 2508 43036 2514
rect 42984 2450 43036 2456
rect 42708 2440 42760 2446
rect 42708 2382 42760 2388
rect 42800 2440 42852 2446
rect 42800 2382 42852 2388
rect 42524 1964 42576 1970
rect 42524 1906 42576 1912
rect 42432 1828 42484 1834
rect 42432 1770 42484 1776
rect 42340 1352 42392 1358
rect 42340 1294 42392 1300
rect 42444 1034 42472 1770
rect 42720 1358 42748 2382
rect 42708 1352 42760 1358
rect 42708 1294 42760 1300
rect 42352 1006 42472 1034
rect 42352 800 42380 1006
rect 42812 800 42840 2382
rect 44188 2202 44540 3238
rect 44640 3052 44692 3058
rect 44640 2994 44692 3000
rect 44652 2650 44680 2994
rect 44640 2644 44692 2650
rect 44640 2586 44692 2592
rect 44188 2150 44210 2202
rect 44262 2150 44274 2202
rect 44326 2150 44338 2202
rect 44390 2150 44402 2202
rect 44454 2150 44466 2202
rect 44518 2150 44540 2202
rect 43720 1896 43772 1902
rect 43720 1838 43772 1844
rect 43260 1828 43312 1834
rect 43260 1770 43312 1776
rect 43272 800 43300 1770
rect 43732 800 43760 1838
rect 43904 1352 43956 1358
rect 43904 1294 43956 1300
rect 43916 1018 43944 1294
rect 44088 1216 44140 1222
rect 44088 1158 44140 1164
rect 44100 1018 44128 1158
rect 44188 1114 44540 2150
rect 44744 2106 44772 4558
rect 44928 3126 44956 5102
rect 45296 5001 45324 5306
rect 45282 4992 45338 5001
rect 45282 4927 45338 4936
rect 45388 4146 45416 5306
rect 45572 5166 45600 5646
rect 47216 5568 47268 5574
rect 47216 5510 47268 5516
rect 47228 5302 47256 5510
rect 47320 5302 47348 6122
rect 47216 5296 47268 5302
rect 47216 5238 47268 5244
rect 47308 5296 47360 5302
rect 47308 5238 47360 5244
rect 45560 5160 45612 5166
rect 45560 5102 45612 5108
rect 47584 5160 47636 5166
rect 47584 5102 47636 5108
rect 45468 5092 45520 5098
rect 45468 5034 45520 5040
rect 45480 4826 45508 5034
rect 45744 5024 45796 5030
rect 45744 4966 45796 4972
rect 45468 4820 45520 4826
rect 45468 4762 45520 4768
rect 45756 4758 45784 4966
rect 45744 4752 45796 4758
rect 45744 4694 45796 4700
rect 46584 4690 46980 4706
rect 46572 4684 46992 4690
rect 46624 4678 46940 4684
rect 46572 4626 46624 4632
rect 46940 4626 46992 4632
rect 46848 4616 46900 4622
rect 46848 4558 46900 4564
rect 45376 4140 45428 4146
rect 45376 4082 45428 4088
rect 46572 4140 46624 4146
rect 46572 4082 46624 4088
rect 46584 4010 46612 4082
rect 46296 4004 46348 4010
rect 46296 3946 46348 3952
rect 46572 4004 46624 4010
rect 46572 3946 46624 3952
rect 45468 3528 45520 3534
rect 45468 3470 45520 3476
rect 45008 3188 45060 3194
rect 45008 3130 45060 3136
rect 44916 3120 44968 3126
rect 44916 3062 44968 3068
rect 45020 3058 45048 3130
rect 45008 3052 45060 3058
rect 45008 2994 45060 3000
rect 45480 2854 45508 3470
rect 46308 3466 46336 3946
rect 46584 3670 46612 3946
rect 46572 3664 46624 3670
rect 46572 3606 46624 3612
rect 46296 3460 46348 3466
rect 46296 3402 46348 3408
rect 46112 3392 46164 3398
rect 46112 3334 46164 3340
rect 46124 3058 46152 3334
rect 46112 3052 46164 3058
rect 46112 2994 46164 3000
rect 45100 2848 45152 2854
rect 45100 2790 45152 2796
rect 45468 2848 45520 2854
rect 45468 2790 45520 2796
rect 45112 2106 45140 2790
rect 45468 2440 45520 2446
rect 45468 2382 45520 2388
rect 44732 2100 44784 2106
rect 44732 2042 44784 2048
rect 45100 2100 45152 2106
rect 45100 2042 45152 2048
rect 45480 1358 45508 2382
rect 46860 2310 46888 4558
rect 47596 3942 47624 5102
rect 48148 3942 48176 6802
rect 50724 5914 50752 7822
rect 59664 7834 59692 8024
rect 59274 7783 59330 7792
rect 59648 7806 59692 7834
rect 62488 7880 62540 7886
rect 62488 7822 62540 7828
rect 63224 7880 63276 7886
rect 63224 7822 63276 7828
rect 59648 7721 59676 7806
rect 59634 7712 59690 7721
rect 59634 7647 59690 7656
rect 61290 7712 61346 7721
rect 61290 7647 61346 7656
rect 61474 7712 61530 7721
rect 61474 7647 61530 7656
rect 58254 7576 58310 7585
rect 58254 7511 58310 7520
rect 58992 7540 59044 7546
rect 57334 7168 57390 7177
rect 57334 7103 57390 7112
rect 55034 6760 55090 6769
rect 55034 6695 55090 6704
rect 51448 6656 51500 6662
rect 51448 6598 51500 6604
rect 52366 6624 52422 6633
rect 51460 5914 51488 6598
rect 52366 6559 52422 6568
rect 52276 6452 52328 6458
rect 52276 6394 52328 6400
rect 50712 5908 50764 5914
rect 50712 5850 50764 5856
rect 51448 5908 51500 5914
rect 51448 5850 51500 5856
rect 49056 5704 49108 5710
rect 49056 5646 49108 5652
rect 50804 5704 50856 5710
rect 50804 5646 50856 5652
rect 51264 5704 51316 5710
rect 51264 5646 51316 5652
rect 51724 5704 51776 5710
rect 51724 5646 51776 5652
rect 48504 5364 48556 5370
rect 48504 5306 48556 5312
rect 48516 5166 48544 5306
rect 48412 5160 48464 5166
rect 48412 5102 48464 5108
rect 48504 5160 48556 5166
rect 48504 5102 48556 5108
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 48136 3936 48188 3942
rect 48136 3878 48188 3884
rect 48136 3664 48188 3670
rect 48136 3606 48188 3612
rect 48148 3466 48176 3606
rect 48044 3460 48096 3466
rect 48044 3402 48096 3408
rect 48136 3460 48188 3466
rect 48136 3402 48188 3408
rect 48056 3346 48084 3402
rect 48056 3318 48176 3346
rect 47676 3052 47728 3058
rect 48044 3052 48096 3058
rect 47728 3012 48044 3040
rect 47676 2994 47728 3000
rect 48044 2994 48096 3000
rect 48148 2990 48176 3318
rect 48136 2984 48188 2990
rect 48136 2926 48188 2932
rect 48424 2582 48452 5102
rect 49068 5030 49096 5646
rect 49056 5024 49108 5030
rect 48502 4992 48558 5001
rect 49056 4966 49108 4972
rect 48502 4927 48558 4936
rect 48412 2576 48464 2582
rect 48412 2518 48464 2524
rect 46940 2440 46992 2446
rect 46940 2382 46992 2388
rect 47400 2440 47452 2446
rect 47400 2382 47452 2388
rect 46848 2304 46900 2310
rect 46848 2246 46900 2252
rect 46952 2106 46980 2382
rect 47032 2304 47084 2310
rect 47032 2246 47084 2252
rect 46940 2100 46992 2106
rect 46940 2042 46992 2048
rect 47044 1970 47072 2246
rect 47032 1964 47084 1970
rect 47032 1906 47084 1912
rect 46020 1896 46072 1902
rect 46020 1838 46072 1844
rect 45192 1352 45244 1358
rect 45192 1294 45244 1300
rect 45468 1352 45520 1358
rect 45468 1294 45520 1300
rect 45100 1284 45152 1290
rect 45100 1226 45152 1232
rect 44640 1216 44692 1222
rect 44640 1158 44692 1164
rect 44188 1062 44210 1114
rect 44262 1062 44274 1114
rect 44326 1062 44338 1114
rect 44390 1062 44402 1114
rect 44454 1062 44466 1114
rect 44518 1062 44540 1114
rect 44188 1040 44540 1062
rect 43904 1012 43956 1018
rect 43904 954 43956 960
rect 44088 1012 44140 1018
rect 44088 954 44140 960
rect 44652 800 44680 1158
rect 45112 800 45140 1226
rect 45204 950 45232 1294
rect 45192 944 45244 950
rect 45192 886 45244 892
rect 46032 800 46060 1838
rect 46480 1284 46532 1290
rect 46480 1226 46532 1232
rect 46492 800 46520 1226
rect 47412 800 47440 2382
rect 48136 2304 48188 2310
rect 48136 2246 48188 2252
rect 47584 2100 47636 2106
rect 47584 2042 47636 2048
rect 47596 1494 47624 2042
rect 47768 1964 47820 1970
rect 47768 1906 47820 1912
rect 47952 1964 48004 1970
rect 47952 1906 48004 1912
rect 47584 1488 47636 1494
rect 47584 1430 47636 1436
rect 47780 1358 47808 1906
rect 47860 1896 47912 1902
rect 47860 1838 47912 1844
rect 47492 1352 47544 1358
rect 47492 1294 47544 1300
rect 47768 1352 47820 1358
rect 47768 1294 47820 1300
rect 47504 882 47532 1294
rect 47492 876 47544 882
rect 47492 818 47544 824
rect 47872 800 47900 1838
rect 47964 1737 47992 1906
rect 47950 1728 48006 1737
rect 47950 1663 48006 1672
rect 48148 1222 48176 2246
rect 48136 1216 48188 1222
rect 48136 1158 48188 1164
rect 48516 950 48544 4927
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 48596 4004 48648 4010
rect 48596 3946 48648 3952
rect 48608 2774 48636 3946
rect 50356 3777 50384 4082
rect 50342 3768 50398 3777
rect 50342 3703 50398 3712
rect 50816 2854 50844 5646
rect 51172 5636 51224 5642
rect 51172 5578 51224 5584
rect 51080 4004 51132 4010
rect 51080 3946 51132 3952
rect 51092 3670 51120 3946
rect 51080 3664 51132 3670
rect 51080 3606 51132 3612
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 50894 3224 50950 3233
rect 51000 3194 51028 3470
rect 51184 3233 51212 5578
rect 51170 3224 51226 3233
rect 50894 3159 50896 3168
rect 50948 3159 50950 3168
rect 50988 3188 51040 3194
rect 50896 3130 50948 3136
rect 51170 3159 51226 3168
rect 50988 3130 51040 3136
rect 50804 2848 50856 2854
rect 50804 2790 50856 2796
rect 48608 2746 48820 2774
rect 48792 2038 48820 2746
rect 49424 2440 49476 2446
rect 49424 2382 49476 2388
rect 50160 2440 50212 2446
rect 50160 2382 50212 2388
rect 49436 2106 49464 2382
rect 49424 2100 49476 2106
rect 49424 2042 49476 2048
rect 48780 2032 48832 2038
rect 48780 1974 48832 1980
rect 48780 1896 48832 1902
rect 48780 1838 48832 1844
rect 48504 944 48556 950
rect 48504 886 48556 892
rect 48792 800 48820 1838
rect 49240 1420 49292 1426
rect 49240 1362 49292 1368
rect 49148 1284 49200 1290
rect 49148 1226 49200 1232
rect 49160 1018 49188 1226
rect 49148 1012 49200 1018
rect 49148 954 49200 960
rect 49252 800 49280 1362
rect 49608 1352 49660 1358
rect 49608 1294 49660 1300
rect 49620 950 49648 1294
rect 49608 944 49660 950
rect 49608 886 49660 892
rect 50172 800 50200 2382
rect 50804 2304 50856 2310
rect 50804 2246 50856 2252
rect 50528 1964 50580 1970
rect 50528 1906 50580 1912
rect 50540 1222 50568 1906
rect 50620 1896 50672 1902
rect 50620 1838 50672 1844
rect 50528 1216 50580 1222
rect 50528 1158 50580 1164
rect 50632 800 50660 1838
rect 50816 1358 50844 2246
rect 51276 1766 51304 5646
rect 51448 4004 51500 4010
rect 51448 3946 51500 3952
rect 51460 3534 51488 3946
rect 51448 3528 51500 3534
rect 51448 3470 51500 3476
rect 51736 3194 51764 5646
rect 51836 4922 52188 5944
rect 52288 5914 52316 6394
rect 52276 5908 52328 5914
rect 52276 5850 52328 5856
rect 51836 4870 51858 4922
rect 51910 4870 51922 4922
rect 51974 4870 51986 4922
rect 52038 4870 52050 4922
rect 52102 4870 52114 4922
rect 52166 4870 52188 4922
rect 51836 3834 52188 4870
rect 52380 3942 52408 6559
rect 53104 6384 53156 6390
rect 53104 6326 53156 6332
rect 53116 6254 53144 6326
rect 53104 6248 53156 6254
rect 53104 6190 53156 6196
rect 53288 6112 53340 6118
rect 53288 6054 53340 6060
rect 53300 5914 53328 6054
rect 53288 5908 53340 5914
rect 53288 5850 53340 5856
rect 52736 5704 52788 5710
rect 52736 5646 52788 5652
rect 52460 5160 52512 5166
rect 52460 5102 52512 5108
rect 52368 3936 52420 3942
rect 52368 3878 52420 3884
rect 51836 3782 51858 3834
rect 51910 3782 51922 3834
rect 51974 3782 51986 3834
rect 52038 3782 52050 3834
rect 52102 3782 52114 3834
rect 52166 3782 52188 3834
rect 51724 3188 51776 3194
rect 51724 3130 51776 3136
rect 51836 2746 52188 3782
rect 52276 3528 52328 3534
rect 52276 3470 52328 3476
rect 51836 2694 51858 2746
rect 51910 2694 51922 2746
rect 51974 2694 51986 2746
rect 52038 2694 52050 2746
rect 52102 2694 52114 2746
rect 52166 2694 52188 2746
rect 51632 2576 51684 2582
rect 51632 2518 51684 2524
rect 51644 2378 51672 2518
rect 51632 2372 51684 2378
rect 51632 2314 51684 2320
rect 51836 2236 52188 2694
rect 51836 2180 51864 2236
rect 51920 2180 51944 2236
rect 52000 2180 52024 2236
rect 52080 2180 52104 2236
rect 52160 2180 52188 2236
rect 51836 2156 52188 2180
rect 51836 2100 51864 2156
rect 51920 2100 51944 2156
rect 52000 2100 52024 2156
rect 52080 2100 52104 2156
rect 52160 2100 52188 2156
rect 51836 2076 52188 2100
rect 51836 2020 51864 2076
rect 51920 2020 51944 2076
rect 52000 2020 52024 2076
rect 52080 2020 52104 2076
rect 52160 2020 52188 2076
rect 51836 1996 52188 2020
rect 51836 1940 51864 1996
rect 51920 1940 51944 1996
rect 52000 1940 52024 1996
rect 52080 1940 52104 1996
rect 52160 1940 52188 1996
rect 51540 1896 51592 1902
rect 51540 1838 51592 1844
rect 51264 1760 51316 1766
rect 51264 1702 51316 1708
rect 50804 1352 50856 1358
rect 50804 1294 50856 1300
rect 51552 800 51580 1838
rect 51836 1658 52188 1940
rect 51836 1606 51858 1658
rect 51910 1606 51922 1658
rect 51974 1606 51986 1658
rect 52038 1606 52050 1658
rect 52102 1606 52114 1658
rect 52166 1606 52188 1658
rect 51724 1284 51776 1290
rect 51724 1226 51776 1232
rect 51736 1018 51764 1226
rect 51836 1040 52188 1606
rect 52288 1358 52316 3470
rect 52472 2650 52500 5102
rect 52748 3398 52776 5646
rect 53746 5536 53802 5545
rect 53746 5471 53802 5480
rect 53760 4554 53788 5471
rect 54188 5466 54540 5944
rect 54188 5414 54210 5466
rect 54262 5414 54274 5466
rect 54326 5414 54338 5466
rect 54390 5414 54402 5466
rect 54454 5414 54466 5466
rect 54518 5414 54540 5466
rect 54188 4588 54540 5414
rect 53748 4548 53800 4554
rect 53748 4490 53800 4496
rect 54188 4532 54216 4588
rect 54272 4532 54296 4588
rect 54352 4532 54376 4588
rect 54432 4532 54456 4588
rect 54512 4532 54540 4588
rect 54188 4508 54540 4532
rect 54188 4452 54216 4508
rect 54272 4452 54296 4508
rect 54352 4452 54376 4508
rect 54432 4452 54456 4508
rect 54512 4452 54540 4508
rect 54188 4428 54540 4452
rect 54188 4378 54216 4428
rect 54272 4378 54296 4428
rect 54352 4378 54376 4428
rect 54432 4378 54456 4428
rect 54512 4378 54540 4428
rect 54188 4326 54210 4378
rect 54272 4372 54274 4378
rect 54454 4372 54456 4378
rect 54262 4348 54274 4372
rect 54326 4348 54338 4372
rect 54390 4348 54402 4372
rect 54454 4348 54466 4372
rect 54272 4326 54274 4348
rect 54454 4326 54456 4348
rect 54518 4326 54540 4378
rect 54188 4292 54216 4326
rect 54272 4292 54296 4326
rect 54352 4292 54376 4326
rect 54432 4292 54456 4326
rect 54512 4292 54540 4326
rect 53380 4072 53432 4078
rect 53380 4014 53432 4020
rect 53104 3664 53156 3670
rect 53104 3606 53156 3612
rect 52736 3392 52788 3398
rect 53012 3392 53064 3398
rect 52736 3334 52788 3340
rect 53010 3360 53012 3369
rect 53064 3360 53066 3369
rect 53010 3295 53066 3304
rect 52460 2644 52512 2650
rect 52460 2586 52512 2592
rect 52644 2440 52696 2446
rect 52644 2382 52696 2388
rect 52656 2106 52684 2382
rect 52644 2100 52696 2106
rect 52644 2042 52696 2048
rect 53116 1970 53144 3606
rect 53392 3369 53420 4014
rect 54024 3936 54076 3942
rect 54024 3878 54076 3884
rect 53378 3360 53434 3369
rect 53378 3295 53434 3304
rect 53656 2440 53708 2446
rect 53656 2382 53708 2388
rect 53104 1964 53156 1970
rect 53104 1906 53156 1912
rect 53380 1896 53432 1902
rect 53380 1838 53432 1844
rect 52276 1352 52328 1358
rect 52276 1294 52328 1300
rect 52368 1284 52420 1290
rect 52368 1226 52420 1232
rect 51724 1012 51776 1018
rect 51724 954 51776 960
rect 52012 870 52132 898
rect 52012 800 52040 870
rect 41984 734 42288 762
rect 42338 0 42394 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44178 0 44234 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47398 0 47454 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 48778 0 48834 800
rect 49238 0 49294 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 50618 0 50674 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 51998 0 52054 800
rect 52104 762 52132 870
rect 52380 762 52408 1226
rect 52920 1216 52972 1222
rect 52920 1158 52972 1164
rect 52932 800 52960 1158
rect 53392 800 53420 1838
rect 53668 1358 53696 2382
rect 54036 1970 54064 3878
rect 54188 3290 54540 4292
rect 55048 4078 55076 6695
rect 56600 6248 56652 6254
rect 56600 6190 56652 6196
rect 56506 5944 56562 5953
rect 56506 5879 56562 5888
rect 55220 5704 55272 5710
rect 55220 5646 55272 5652
rect 55956 5704 56008 5710
rect 55956 5646 56008 5652
rect 55036 4072 55088 4078
rect 55036 4014 55088 4020
rect 54852 3936 54904 3942
rect 54852 3878 54904 3884
rect 54188 3238 54210 3290
rect 54262 3238 54274 3290
rect 54326 3238 54338 3290
rect 54390 3238 54402 3290
rect 54454 3238 54466 3290
rect 54518 3238 54540 3290
rect 54188 2202 54540 3238
rect 54188 2150 54210 2202
rect 54262 2150 54274 2202
rect 54326 2150 54338 2202
rect 54390 2150 54402 2202
rect 54454 2150 54466 2202
rect 54518 2150 54540 2202
rect 54024 1964 54076 1970
rect 54024 1906 54076 1912
rect 53656 1352 53708 1358
rect 53656 1294 53708 1300
rect 54188 1114 54540 2150
rect 54576 1896 54628 1902
rect 54576 1838 54628 1844
rect 54188 1062 54210 1114
rect 54262 1062 54274 1114
rect 54326 1062 54338 1114
rect 54390 1062 54402 1114
rect 54454 1062 54466 1114
rect 54518 1062 54540 1114
rect 54188 1040 54540 1062
rect 54312 870 54432 898
rect 54312 800 54340 870
rect 52104 734 52408 762
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 53838 0 53894 800
rect 54298 0 54354 800
rect 54404 762 54432 870
rect 54588 762 54616 1838
rect 54864 1358 54892 3878
rect 55232 1834 55260 5646
rect 55588 2440 55640 2446
rect 55588 2382 55640 2388
rect 55600 2106 55628 2382
rect 55772 2304 55824 2310
rect 55772 2246 55824 2252
rect 55588 2100 55640 2106
rect 55588 2042 55640 2048
rect 55784 1970 55812 2246
rect 55772 1964 55824 1970
rect 55772 1906 55824 1912
rect 55220 1828 55272 1834
rect 55220 1770 55272 1776
rect 55968 1494 55996 5646
rect 56520 4078 56548 5879
rect 56612 5710 56640 6190
rect 57348 5778 57376 7103
rect 57336 5772 57388 5778
rect 57336 5714 57388 5720
rect 56600 5704 56652 5710
rect 56600 5646 56652 5652
rect 56692 5704 56744 5710
rect 56692 5646 56744 5652
rect 56508 4072 56560 4078
rect 56508 4014 56560 4020
rect 56704 2514 56732 5646
rect 58268 4078 58296 7511
rect 58992 7482 59044 7488
rect 58900 7336 58952 7342
rect 58900 7278 58952 7284
rect 58912 5030 58940 7278
rect 58900 5024 58952 5030
rect 58900 4966 58952 4972
rect 58256 4072 58308 4078
rect 58256 4014 58308 4020
rect 57428 4004 57480 4010
rect 57428 3946 57480 3952
rect 56692 2508 56744 2514
rect 56692 2450 56744 2456
rect 57440 2446 57468 3946
rect 57612 3936 57664 3942
rect 57612 3878 57664 3884
rect 58440 3936 58492 3942
rect 58440 3878 58492 3884
rect 57624 3534 57652 3878
rect 58452 3670 58480 3878
rect 58440 3664 58492 3670
rect 58440 3606 58492 3612
rect 57796 3596 57848 3602
rect 57796 3538 57848 3544
rect 57612 3528 57664 3534
rect 57612 3470 57664 3476
rect 57808 3194 57836 3538
rect 58716 3460 58768 3466
rect 58716 3402 58768 3408
rect 58900 3460 58952 3466
rect 58900 3402 58952 3408
rect 58728 3233 58756 3402
rect 58714 3224 58770 3233
rect 57796 3188 57848 3194
rect 58714 3159 58770 3168
rect 57796 3130 57848 3136
rect 57520 2508 57572 2514
rect 57520 2450 57572 2456
rect 56324 2440 56376 2446
rect 56324 2382 56376 2388
rect 57428 2440 57480 2446
rect 57428 2382 57480 2388
rect 56140 1896 56192 1902
rect 56140 1838 56192 1844
rect 55956 1488 56008 1494
rect 55956 1430 56008 1436
rect 54852 1352 54904 1358
rect 54852 1294 54904 1300
rect 54760 1284 54812 1290
rect 54760 1226 54812 1232
rect 54772 800 54800 1226
rect 55680 1216 55732 1222
rect 55680 1158 55732 1164
rect 55692 800 55720 1158
rect 56152 800 56180 1838
rect 56336 1358 56364 2382
rect 57060 1964 57112 1970
rect 57060 1906 57112 1912
rect 56324 1352 56376 1358
rect 56324 1294 56376 1300
rect 57072 800 57100 1906
rect 57336 1216 57388 1222
rect 57336 1158 57388 1164
rect 57348 1018 57376 1158
rect 57336 1012 57388 1018
rect 57336 954 57388 960
rect 57532 800 57560 2450
rect 58532 2440 58584 2446
rect 58532 2382 58584 2388
rect 58440 1760 58492 1766
rect 58440 1702 58492 1708
rect 58452 1426 58480 1702
rect 58440 1420 58492 1426
rect 58440 1362 58492 1368
rect 58544 1306 58572 2382
rect 58452 1278 58572 1306
rect 58452 800 58480 1278
rect 58912 800 58940 3402
rect 59004 3194 59032 7482
rect 61304 7449 61332 7647
rect 61290 7440 61346 7449
rect 60004 7404 60056 7410
rect 61290 7375 61346 7384
rect 60004 7346 60056 7352
rect 59084 7268 59136 7274
rect 59084 7210 59136 7216
rect 59096 5370 59124 7210
rect 59544 7200 59596 7206
rect 59544 7142 59596 7148
rect 59268 7132 59320 7138
rect 59268 7074 59320 7080
rect 59176 5908 59228 5914
rect 59176 5850 59228 5856
rect 59084 5364 59136 5370
rect 59084 5306 59136 5312
rect 59188 5030 59216 5850
rect 59176 5024 59228 5030
rect 59176 4966 59228 4972
rect 59188 4486 59216 4966
rect 59280 4758 59308 7074
rect 59360 6996 59412 7002
rect 59360 6938 59412 6944
rect 59268 4752 59320 4758
rect 59268 4694 59320 4700
rect 59372 4690 59400 6938
rect 59360 4684 59412 4690
rect 59360 4626 59412 4632
rect 59556 4554 59584 7142
rect 59728 7064 59780 7070
rect 59728 7006 59780 7012
rect 59740 5914 59768 7006
rect 59728 5908 59780 5914
rect 59728 5850 59780 5856
rect 60016 4622 60044 7346
rect 61200 6928 61252 6934
rect 61200 6870 61252 6876
rect 60740 5908 60792 5914
rect 60740 5850 60792 5856
rect 60844 5902 61148 5930
rect 61212 5914 61240 6870
rect 61488 6118 61516 7647
rect 61476 6112 61528 6118
rect 61476 6054 61528 6060
rect 60280 5160 60332 5166
rect 60278 5128 60280 5137
rect 60332 5128 60334 5137
rect 60278 5063 60334 5072
rect 60752 5030 60780 5850
rect 60844 5778 60872 5902
rect 61120 5794 61148 5902
rect 61200 5908 61252 5914
rect 61200 5850 61252 5856
rect 61292 5908 61344 5914
rect 61292 5850 61344 5856
rect 61304 5794 61332 5850
rect 60832 5772 60884 5778
rect 61120 5766 61332 5794
rect 60832 5714 60884 5720
rect 61752 5296 61804 5302
rect 61750 5264 61752 5273
rect 61804 5264 61806 5273
rect 61750 5199 61806 5208
rect 61108 5092 61160 5098
rect 61108 5034 61160 5040
rect 60740 5024 60792 5030
rect 60462 4992 60518 5001
rect 61120 5001 61148 5034
rect 60740 4966 60792 4972
rect 61106 4992 61162 5001
rect 60462 4927 60518 4936
rect 60476 4826 60504 4927
rect 60464 4820 60516 4826
rect 60464 4762 60516 4768
rect 60004 4616 60056 4622
rect 60004 4558 60056 4564
rect 60648 4616 60700 4622
rect 60648 4558 60700 4564
rect 59544 4548 59596 4554
rect 59544 4490 59596 4496
rect 59176 4480 59228 4486
rect 59176 4422 59228 4428
rect 59360 4480 59412 4486
rect 59360 4422 59412 4428
rect 59188 4078 59216 4422
rect 59372 4282 59400 4422
rect 59360 4276 59412 4282
rect 59360 4218 59412 4224
rect 60556 4276 60608 4282
rect 60556 4218 60608 4224
rect 59176 4072 59228 4078
rect 59176 4014 59228 4020
rect 59188 3398 59216 4014
rect 60568 3398 60596 4218
rect 60660 4146 60688 4558
rect 60752 4554 60780 4966
rect 61106 4927 61162 4936
rect 61836 4922 62188 5972
rect 62304 5568 62356 5574
rect 62304 5510 62356 5516
rect 62316 5302 62344 5510
rect 62304 5296 62356 5302
rect 62396 5296 62448 5302
rect 62304 5238 62356 5244
rect 62394 5264 62396 5273
rect 62448 5264 62450 5273
rect 61836 4870 61858 4922
rect 61910 4870 61922 4922
rect 61974 4870 61986 4922
rect 62038 4870 62050 4922
rect 62102 4870 62114 4922
rect 62166 4870 62188 4922
rect 61200 4752 61252 4758
rect 61200 4694 61252 4700
rect 60740 4548 60792 4554
rect 60740 4490 60792 4496
rect 60752 4282 60780 4490
rect 60832 4480 60884 4486
rect 60832 4422 60884 4428
rect 60924 4480 60976 4486
rect 60924 4422 60976 4428
rect 60844 4282 60872 4422
rect 60740 4276 60792 4282
rect 60740 4218 60792 4224
rect 60832 4276 60884 4282
rect 60832 4218 60884 4224
rect 60936 4214 60964 4422
rect 60924 4208 60976 4214
rect 61212 4185 61240 4694
rect 61476 4548 61528 4554
rect 61476 4490 61528 4496
rect 60924 4150 60976 4156
rect 61198 4176 61254 4185
rect 60648 4140 60700 4146
rect 61198 4111 61254 4120
rect 60648 4082 60700 4088
rect 60648 3732 60700 3738
rect 60648 3674 60700 3680
rect 60660 3398 60688 3674
rect 61488 3534 61516 4490
rect 61660 4004 61712 4010
rect 61660 3946 61712 3952
rect 61568 3664 61620 3670
rect 61568 3606 61620 3612
rect 61476 3528 61528 3534
rect 61476 3470 61528 3476
rect 59176 3392 59228 3398
rect 59176 3334 59228 3340
rect 60556 3392 60608 3398
rect 60556 3334 60608 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 59188 3210 59216 3334
rect 59096 3194 59216 3210
rect 58992 3188 59044 3194
rect 58992 3130 59044 3136
rect 59084 3188 59216 3194
rect 59136 3182 59216 3188
rect 59084 3130 59136 3136
rect 59096 2514 59124 3130
rect 60568 3126 60596 3334
rect 59176 3120 59228 3126
rect 59176 3062 59228 3068
rect 60556 3120 60608 3126
rect 60556 3062 60608 3068
rect 59188 2854 59216 3062
rect 59268 3052 59320 3058
rect 59268 2994 59320 3000
rect 59636 3052 59688 3058
rect 59636 2994 59688 3000
rect 59176 2848 59228 2854
rect 59176 2790 59228 2796
rect 59084 2508 59136 2514
rect 59084 2450 59136 2456
rect 59096 2106 59124 2450
rect 59176 2304 59228 2310
rect 59176 2246 59228 2252
rect 59084 2100 59136 2106
rect 59084 2042 59136 2048
rect 59096 1562 59124 2042
rect 59188 1562 59216 2246
rect 59084 1556 59136 1562
rect 59084 1498 59136 1504
rect 59176 1556 59228 1562
rect 59176 1498 59228 1504
rect 59280 1358 59308 2994
rect 59648 2106 59676 2994
rect 60568 2514 60596 3062
rect 61580 3058 61608 3606
rect 61568 3052 61620 3058
rect 61568 2994 61620 3000
rect 61672 2514 61700 3946
rect 61836 3834 62188 4870
rect 62316 4826 62344 5238
rect 62394 5199 62450 5208
rect 62304 4820 62356 4826
rect 62304 4762 62356 4768
rect 62316 4078 62344 4762
rect 62304 4072 62356 4078
rect 62304 4014 62356 4020
rect 61836 3782 61858 3834
rect 61910 3782 61922 3834
rect 61974 3782 61986 3834
rect 62038 3782 62050 3834
rect 62102 3782 62114 3834
rect 62166 3782 62188 3834
rect 61836 2746 62188 3782
rect 62316 3670 62344 4014
rect 62304 3664 62356 3670
rect 62304 3606 62356 3612
rect 62316 3126 62344 3606
rect 62396 3392 62448 3398
rect 62396 3334 62448 3340
rect 62408 3233 62436 3334
rect 62394 3224 62450 3233
rect 62500 3194 62528 7822
rect 63236 7698 63264 7822
rect 63408 7812 63460 7818
rect 63408 7754 63460 7760
rect 62960 7670 63264 7698
rect 62670 7304 62726 7313
rect 62670 7239 62726 7248
rect 62578 7032 62634 7041
rect 62578 6967 62634 6976
rect 62592 3466 62620 6967
rect 62684 4026 62712 7239
rect 62856 6724 62908 6730
rect 62856 6666 62908 6672
rect 62868 6390 62896 6666
rect 62764 6384 62816 6390
rect 62764 6326 62816 6332
rect 62856 6384 62908 6390
rect 62856 6326 62908 6332
rect 62776 6118 62804 6326
rect 62764 6112 62816 6118
rect 62764 6054 62816 6060
rect 62854 6080 62910 6089
rect 62854 6015 62910 6024
rect 62868 5642 62896 6015
rect 62856 5636 62908 5642
rect 62856 5578 62908 5584
rect 62764 5160 62816 5166
rect 62764 5102 62816 5108
rect 62776 4486 62804 5102
rect 62764 4480 62816 4486
rect 62764 4422 62816 4428
rect 62684 3998 62804 4026
rect 62672 3936 62724 3942
rect 62672 3878 62724 3884
rect 62580 3460 62632 3466
rect 62580 3402 62632 3408
rect 62394 3159 62450 3168
rect 62488 3188 62540 3194
rect 62488 3130 62540 3136
rect 62304 3120 62356 3126
rect 62356 3080 62436 3108
rect 62304 3062 62356 3068
rect 61836 2694 61858 2746
rect 61910 2694 61922 2746
rect 61974 2694 61986 2746
rect 62038 2694 62050 2746
rect 62102 2694 62114 2746
rect 62166 2694 62188 2746
rect 60556 2508 60608 2514
rect 60556 2450 60608 2456
rect 61660 2508 61712 2514
rect 61660 2450 61712 2456
rect 60096 2372 60148 2378
rect 60096 2314 60148 2320
rect 60004 2304 60056 2310
rect 60004 2246 60056 2252
rect 59636 2100 59688 2106
rect 59636 2042 59688 2048
rect 60016 1970 60044 2246
rect 60108 1970 60136 2314
rect 60568 2106 60596 2450
rect 61384 2440 61436 2446
rect 61384 2382 61436 2388
rect 61016 2304 61068 2310
rect 61016 2246 61068 2252
rect 60556 2100 60608 2106
rect 60556 2042 60608 2048
rect 60004 1964 60056 1970
rect 60004 1906 60056 1912
rect 60096 1964 60148 1970
rect 60096 1906 60148 1912
rect 59820 1896 59872 1902
rect 59820 1838 59872 1844
rect 59268 1352 59320 1358
rect 59268 1294 59320 1300
rect 59832 800 59860 1838
rect 60568 1494 60596 2042
rect 61028 1902 61056 2246
rect 61396 2106 61424 2382
rect 61660 2304 61712 2310
rect 61660 2246 61712 2252
rect 61384 2100 61436 2106
rect 61384 2042 61436 2048
rect 61016 1896 61068 1902
rect 61016 1838 61068 1844
rect 60556 1488 60608 1494
rect 60556 1430 60608 1436
rect 61200 1352 61252 1358
rect 61200 1294 61252 1300
rect 60280 1012 60332 1018
rect 60280 954 60332 960
rect 60292 800 60320 954
rect 61212 800 61240 1294
rect 61672 800 61700 2246
rect 61836 2236 62188 2694
rect 62304 2440 62356 2446
rect 62304 2382 62356 2388
rect 61836 2180 61864 2236
rect 61920 2180 61944 2236
rect 62000 2180 62024 2236
rect 62080 2180 62104 2236
rect 62160 2180 62188 2236
rect 61836 2156 62188 2180
rect 61836 2100 61864 2156
rect 61920 2100 61944 2156
rect 62000 2100 62024 2156
rect 62080 2100 62104 2156
rect 62160 2100 62188 2156
rect 61836 2076 62188 2100
rect 61836 2020 61864 2076
rect 61920 2020 61944 2076
rect 62000 2020 62024 2076
rect 62080 2020 62104 2076
rect 62160 2020 62188 2076
rect 61836 1996 62188 2020
rect 61836 1940 61864 1996
rect 61920 1940 61944 1996
rect 62000 1940 62024 1996
rect 62080 1940 62104 1996
rect 62160 1940 62188 1996
rect 61836 1658 62188 1940
rect 61836 1606 61858 1658
rect 61910 1606 61922 1658
rect 61974 1606 61986 1658
rect 62038 1606 62050 1658
rect 62102 1606 62114 1658
rect 62166 1606 62188 1658
rect 61836 1040 62188 1606
rect 62316 1358 62344 2382
rect 62408 2310 62436 3080
rect 62684 3058 62712 3878
rect 62672 3052 62724 3058
rect 62672 2994 62724 3000
rect 62776 2854 62804 3998
rect 62764 2848 62816 2854
rect 62764 2790 62816 2796
rect 62672 2576 62724 2582
rect 62672 2518 62724 2524
rect 62396 2304 62448 2310
rect 62396 2246 62448 2252
rect 62580 2304 62632 2310
rect 62580 2246 62632 2252
rect 62408 2038 62436 2246
rect 62592 2038 62620 2246
rect 62684 2038 62712 2518
rect 62396 2032 62448 2038
rect 62396 1974 62448 1980
rect 62580 2032 62632 2038
rect 62580 1974 62632 1980
rect 62672 2032 62724 2038
rect 62672 1974 62724 1980
rect 62408 1494 62436 1974
rect 62960 1970 62988 7670
rect 63132 2304 63184 2310
rect 63132 2246 63184 2252
rect 63144 1970 63172 2246
rect 62948 1964 63000 1970
rect 62948 1906 63000 1912
rect 63132 1964 63184 1970
rect 63132 1906 63184 1912
rect 63224 1896 63276 1902
rect 63224 1838 63276 1844
rect 62396 1488 62448 1494
rect 62396 1430 62448 1436
rect 62304 1352 62356 1358
rect 62304 1294 62356 1300
rect 62580 1352 62632 1358
rect 62580 1294 62632 1300
rect 62592 800 62620 1294
rect 63236 1034 63264 1838
rect 63420 1766 63448 7754
rect 63512 6934 63540 9823
rect 63500 6928 63552 6934
rect 63500 6870 63552 6876
rect 63604 6089 63632 10220
rect 63696 7614 63724 12378
rect 63684 7608 63736 7614
rect 63684 7550 63736 7556
rect 63590 6080 63646 6089
rect 63590 6015 63646 6024
rect 63500 5908 63552 5914
rect 63500 5850 63552 5856
rect 63592 5908 63644 5914
rect 63592 5850 63644 5856
rect 63512 5574 63540 5850
rect 63500 5568 63552 5574
rect 63500 5510 63552 5516
rect 63604 5030 63632 5850
rect 63788 5098 63816 42774
rect 63880 41313 63908 74530
rect 64144 73976 64196 73982
rect 64144 73918 64196 73924
rect 63960 63640 64012 63646
rect 63960 63582 64012 63588
rect 63972 62082 64000 63582
rect 63960 62076 64012 62082
rect 63960 62018 64012 62024
rect 63960 61328 64012 61334
rect 63960 61270 64012 61276
rect 63972 55282 64000 61270
rect 63960 55276 64012 55282
rect 63960 55218 64012 55224
rect 64052 54800 64104 54806
rect 64052 54742 64104 54748
rect 64064 43450 64092 54742
rect 64052 43444 64104 43450
rect 64052 43386 64104 43392
rect 63866 41304 63922 41313
rect 63866 41239 63922 41248
rect 63960 40996 64012 41002
rect 63960 40938 64012 40944
rect 63868 38684 63920 38690
rect 63868 38626 63920 38632
rect 63880 5302 63908 38626
rect 63972 17218 64000 40938
rect 64052 38752 64104 38758
rect 64052 38694 64104 38700
rect 64064 17354 64092 38694
rect 64156 17474 64184 73918
rect 65628 71602 65656 78678
rect 65708 72208 65760 72214
rect 65708 72150 65760 72156
rect 65616 71596 65668 71602
rect 65616 71538 65668 71544
rect 65616 70032 65668 70038
rect 65616 69974 65668 69980
rect 64788 67652 64840 67658
rect 64788 67594 64840 67600
rect 64696 52692 64748 52698
rect 64696 52634 64748 52640
rect 64328 48816 64380 48822
rect 64328 48758 64380 48764
rect 64236 44736 64288 44742
rect 64236 44678 64288 44684
rect 64248 31754 64276 44678
rect 64236 31748 64288 31754
rect 64236 31690 64288 31696
rect 64236 31544 64288 31550
rect 64236 31486 64288 31492
rect 64144 17468 64196 17474
rect 64144 17410 64196 17416
rect 64064 17326 64184 17354
rect 63972 17190 64092 17218
rect 63960 12028 64012 12034
rect 63960 11970 64012 11976
rect 63972 7070 64000 11970
rect 64064 7750 64092 17190
rect 64052 7744 64104 7750
rect 64052 7686 64104 7692
rect 64156 7682 64184 17326
rect 64248 7954 64276 31486
rect 64236 7948 64288 7954
rect 64236 7890 64288 7896
rect 64144 7676 64196 7682
rect 64144 7618 64196 7624
rect 63960 7064 64012 7070
rect 63960 7006 64012 7012
rect 64236 6792 64288 6798
rect 64236 6734 64288 6740
rect 64248 6118 64276 6734
rect 64340 6497 64368 48758
rect 64420 47728 64472 47734
rect 64420 47670 64472 47676
rect 64432 31634 64460 47670
rect 64604 43852 64656 43858
rect 64604 43794 64656 43800
rect 64512 36576 64564 36582
rect 64512 36518 64564 36524
rect 64524 31754 64552 36518
rect 64616 31772 64644 43794
rect 64708 40050 64736 52634
rect 64696 40044 64748 40050
rect 64696 39986 64748 39992
rect 64696 33992 64748 33998
rect 64696 33934 64748 33940
rect 64604 31766 64656 31772
rect 64512 31748 64564 31754
rect 64604 31708 64656 31714
rect 64512 31690 64564 31696
rect 64432 31606 64644 31634
rect 64420 31544 64472 31550
rect 64420 31486 64472 31492
rect 64512 31544 64564 31550
rect 64512 31486 64564 31492
rect 64432 30394 64460 31486
rect 64420 30388 64472 30394
rect 64420 30330 64472 30336
rect 64420 27940 64472 27946
rect 64420 27882 64472 27888
rect 64432 22166 64460 27882
rect 64524 22370 64552 31486
rect 64616 25498 64644 31606
rect 64604 25492 64656 25498
rect 64604 25434 64656 25440
rect 64604 25288 64656 25294
rect 64604 25230 64656 25236
rect 64616 22370 64644 25230
rect 64512 22364 64564 22370
rect 64512 22306 64564 22312
rect 64604 22364 64656 22370
rect 64604 22306 64656 22312
rect 64420 22160 64472 22166
rect 64420 22102 64472 22108
rect 64512 22160 64564 22166
rect 64512 22102 64564 22108
rect 64420 22024 64472 22030
rect 64420 21966 64472 21972
rect 64326 6488 64382 6497
rect 64432 6458 64460 21966
rect 64524 6594 64552 22102
rect 64604 22092 64656 22098
rect 64604 22034 64656 22040
rect 64616 17610 64644 22034
rect 64604 17604 64656 17610
rect 64604 17546 64656 17552
rect 64604 17468 64656 17474
rect 64604 17410 64656 17416
rect 64616 11898 64644 17410
rect 64604 11892 64656 11898
rect 64604 11834 64656 11840
rect 64602 11792 64658 11801
rect 64602 11727 64658 11736
rect 64616 7721 64644 11727
rect 64602 7712 64658 7721
rect 64602 7647 64658 7656
rect 64604 6860 64656 6866
rect 64604 6802 64656 6808
rect 64512 6588 64564 6594
rect 64512 6530 64564 6536
rect 64326 6423 64382 6432
rect 64420 6452 64472 6458
rect 64420 6394 64472 6400
rect 64052 6112 64104 6118
rect 64052 6054 64104 6060
rect 64236 6112 64288 6118
rect 64236 6054 64288 6060
rect 64064 5778 64092 6054
rect 64052 5772 64104 5778
rect 64052 5714 64104 5720
rect 64188 5466 64540 5972
rect 64188 5414 64210 5466
rect 64262 5414 64274 5466
rect 64326 5414 64338 5466
rect 64390 5414 64402 5466
rect 64454 5414 64466 5466
rect 64518 5414 64540 5466
rect 63868 5296 63920 5302
rect 63868 5238 63920 5244
rect 63776 5092 63828 5098
rect 63776 5034 63828 5040
rect 63592 5024 63644 5030
rect 63592 4966 63644 4972
rect 63604 4758 63632 4966
rect 63592 4752 63644 4758
rect 63592 4694 63644 4700
rect 63960 4752 64012 4758
rect 63960 4694 64012 4700
rect 63972 4214 64000 4694
rect 64188 4588 64540 5414
rect 64188 4532 64216 4588
rect 64272 4532 64296 4588
rect 64352 4532 64376 4588
rect 64432 4532 64456 4588
rect 64512 4532 64540 4588
rect 64188 4508 64540 4532
rect 64188 4452 64216 4508
rect 64272 4452 64296 4508
rect 64352 4452 64376 4508
rect 64432 4452 64456 4508
rect 64512 4452 64540 4508
rect 64188 4428 64540 4452
rect 64188 4378 64216 4428
rect 64272 4378 64296 4428
rect 64352 4378 64376 4428
rect 64432 4378 64456 4428
rect 64512 4378 64540 4428
rect 64188 4326 64210 4378
rect 64272 4372 64274 4378
rect 64454 4372 64456 4378
rect 64262 4348 64274 4372
rect 64326 4348 64338 4372
rect 64390 4348 64402 4372
rect 64454 4348 64466 4372
rect 64272 4326 64274 4348
rect 64454 4326 64456 4348
rect 64518 4326 64540 4378
rect 64188 4292 64216 4326
rect 64272 4292 64296 4326
rect 64352 4292 64376 4326
rect 64432 4292 64456 4326
rect 64512 4292 64540 4326
rect 63960 4208 64012 4214
rect 63682 4176 63738 4185
rect 63960 4150 64012 4156
rect 63682 4111 63738 4120
rect 63500 3664 63552 3670
rect 63500 3606 63552 3612
rect 63512 3194 63540 3606
rect 63500 3188 63552 3194
rect 63500 3130 63552 3136
rect 63512 2650 63540 3130
rect 63592 3120 63644 3126
rect 63592 3062 63644 3068
rect 63500 2644 63552 2650
rect 63500 2586 63552 2592
rect 63512 1970 63540 2586
rect 63500 1964 63552 1970
rect 63500 1906 63552 1912
rect 63408 1760 63460 1766
rect 63408 1702 63460 1708
rect 63512 1494 63540 1906
rect 63500 1488 63552 1494
rect 63500 1430 63552 1436
rect 63604 1340 63632 3062
rect 63696 1970 63724 4111
rect 63868 4004 63920 4010
rect 63868 3946 63920 3952
rect 63880 2990 63908 3946
rect 63972 3670 64000 4150
rect 63960 3664 64012 3670
rect 63960 3606 64012 3612
rect 64188 3290 64540 4292
rect 64188 3238 64210 3290
rect 64262 3238 64274 3290
rect 64326 3238 64338 3290
rect 64390 3238 64402 3290
rect 64454 3238 64466 3290
rect 64518 3238 64540 3290
rect 63868 2984 63920 2990
rect 63868 2926 63920 2932
rect 63960 2984 64012 2990
rect 63960 2926 64012 2932
rect 63776 2576 63828 2582
rect 63776 2518 63828 2524
rect 63684 1964 63736 1970
rect 63684 1906 63736 1912
rect 63788 1834 63816 2518
rect 63776 1828 63828 1834
rect 63776 1770 63828 1776
rect 63684 1352 63736 1358
rect 63604 1312 63684 1340
rect 63684 1294 63736 1300
rect 63052 1006 63264 1034
rect 63052 800 63080 1006
rect 63972 800 64000 2926
rect 64188 2202 64540 3238
rect 64616 2310 64644 6802
rect 64708 5710 64736 33934
rect 64800 12034 64828 67594
rect 65432 67584 65484 67590
rect 65432 67526 65484 67532
rect 65340 65680 65392 65686
rect 65340 65622 65392 65628
rect 65248 62076 65300 62082
rect 65248 62018 65300 62024
rect 65156 59152 65208 59158
rect 65156 59094 65208 59100
rect 65064 56976 65116 56982
rect 65064 56918 65116 56924
rect 64972 55276 65024 55282
rect 64972 55218 65024 55224
rect 64880 50448 64932 50454
rect 64880 50390 64932 50396
rect 64892 26586 64920 50390
rect 64984 32026 65012 55218
rect 65076 40186 65104 56918
rect 65064 40180 65116 40186
rect 65064 40122 65116 40128
rect 65168 40032 65196 59094
rect 65076 40004 65196 40032
rect 64972 32020 65024 32026
rect 64972 31962 65024 31968
rect 65076 30938 65104 40004
rect 65260 39930 65288 62018
rect 65168 39902 65288 39930
rect 65168 33114 65196 39902
rect 65352 39794 65380 65622
rect 65260 39766 65380 39794
rect 65260 34202 65288 39766
rect 65444 39658 65472 67526
rect 65524 47524 65576 47530
rect 65524 47466 65576 47472
rect 65536 43654 65564 47466
rect 65524 43648 65576 43654
rect 65524 43590 65576 43596
rect 65524 43444 65576 43450
rect 65524 43386 65576 43392
rect 65536 40594 65564 43386
rect 65524 40588 65576 40594
rect 65524 40530 65576 40536
rect 65524 40044 65576 40050
rect 65524 39986 65576 39992
rect 65352 39630 65472 39658
rect 65352 34746 65380 39630
rect 65536 39522 65564 39986
rect 65444 39494 65564 39522
rect 65444 36258 65472 39494
rect 65628 39386 65656 69974
rect 65720 55214 65748 72150
rect 66168 71664 66220 71670
rect 66168 71606 66220 71612
rect 65720 55186 65840 55214
rect 65708 47048 65760 47054
rect 65706 47016 65708 47025
rect 65760 47016 65762 47025
rect 65706 46951 65762 46960
rect 65812 46866 65840 55186
rect 66076 47116 66128 47122
rect 66076 47058 66128 47064
rect 65984 47048 66036 47054
rect 65982 47016 65984 47025
rect 66036 47016 66038 47025
rect 65982 46951 66038 46960
rect 65536 39358 65656 39386
rect 65720 46838 65840 46866
rect 65536 36378 65564 39358
rect 65720 39250 65748 46838
rect 65800 45960 65852 45966
rect 65800 45902 65852 45908
rect 65628 39222 65748 39250
rect 65628 38010 65656 39222
rect 65706 38584 65762 38593
rect 65706 38519 65708 38528
rect 65760 38519 65762 38528
rect 65708 38490 65760 38496
rect 65616 38004 65668 38010
rect 65616 37946 65668 37952
rect 65524 36372 65576 36378
rect 65524 36314 65576 36320
rect 65444 36230 65656 36258
rect 65432 36168 65484 36174
rect 65432 36110 65484 36116
rect 65524 36168 65576 36174
rect 65524 36110 65576 36116
rect 65444 35222 65472 36110
rect 65432 35216 65484 35222
rect 65432 35158 65484 35164
rect 65432 35080 65484 35086
rect 65432 35022 65484 35028
rect 65444 34785 65472 35022
rect 65430 34776 65486 34785
rect 65340 34740 65392 34746
rect 65430 34711 65486 34720
rect 65340 34682 65392 34688
rect 65340 34604 65392 34610
rect 65340 34546 65392 34552
rect 65248 34196 65300 34202
rect 65248 34138 65300 34144
rect 65156 33108 65208 33114
rect 65156 33050 65208 33056
rect 65352 31754 65380 34546
rect 65536 31754 65564 36110
rect 65260 31726 65380 31754
rect 65444 31726 65564 31754
rect 65064 30932 65116 30938
rect 65064 30874 65116 30880
rect 65156 30864 65208 30870
rect 65156 30806 65208 30812
rect 64972 30388 65024 30394
rect 64972 30330 65024 30336
rect 64880 26580 64932 26586
rect 64880 26522 64932 26528
rect 64880 24336 64932 24342
rect 64880 24278 64932 24284
rect 64892 22574 64920 24278
rect 64880 22568 64932 22574
rect 64880 22510 64932 22516
rect 64880 22364 64932 22370
rect 64880 22306 64932 22312
rect 64892 22030 64920 22306
rect 64880 22024 64932 22030
rect 64880 21966 64932 21972
rect 64880 19304 64932 19310
rect 64880 19246 64932 19252
rect 64892 18086 64920 19246
rect 64880 18080 64932 18086
rect 64880 18022 64932 18028
rect 64880 12504 64932 12510
rect 64880 12446 64932 12452
rect 64788 12028 64840 12034
rect 64788 11970 64840 11976
rect 64788 11892 64840 11898
rect 64788 11834 64840 11840
rect 64800 7546 64828 11834
rect 64788 7540 64840 7546
rect 64788 7482 64840 7488
rect 64800 5914 64828 7482
rect 64892 6254 64920 12446
rect 64880 6248 64932 6254
rect 64880 6190 64932 6196
rect 64788 5908 64840 5914
rect 64788 5850 64840 5856
rect 64696 5704 64748 5710
rect 64696 5646 64748 5652
rect 64788 5704 64840 5710
rect 64788 5646 64840 5652
rect 64800 3738 64828 5646
rect 64984 4162 65012 30330
rect 65168 28694 65196 30806
rect 65156 28688 65208 28694
rect 65156 28630 65208 28636
rect 65168 26790 65196 28630
rect 65156 26784 65208 26790
rect 65156 26726 65208 26732
rect 65064 17604 65116 17610
rect 65064 17546 65116 17552
rect 65076 12442 65104 17546
rect 65064 12436 65116 12442
rect 65064 12378 65116 12384
rect 65064 11892 65116 11898
rect 65064 11834 65116 11840
rect 65076 4554 65104 11834
rect 65168 7138 65196 26726
rect 65260 23798 65288 31726
rect 65444 28914 65472 31726
rect 65352 28886 65472 28914
rect 65352 28218 65380 28886
rect 65628 28778 65656 36230
rect 65708 35692 65760 35698
rect 65708 35634 65760 35640
rect 65444 28750 65656 28778
rect 65340 28212 65392 28218
rect 65340 28154 65392 28160
rect 65444 27606 65472 28750
rect 65720 28642 65748 35634
rect 65536 28614 65748 28642
rect 65536 28422 65564 28614
rect 65708 28484 65760 28490
rect 65708 28426 65760 28432
rect 65524 28416 65576 28422
rect 65524 28358 65576 28364
rect 65432 27600 65484 27606
rect 65432 27542 65484 27548
rect 65432 25288 65484 25294
rect 65432 25230 65484 25236
rect 65444 24614 65472 25230
rect 65432 24608 65484 24614
rect 65432 24550 65484 24556
rect 65248 23792 65300 23798
rect 65248 23734 65300 23740
rect 65340 23656 65392 23662
rect 65340 23598 65392 23604
rect 65352 22982 65380 23598
rect 65340 22976 65392 22982
rect 65340 22918 65392 22924
rect 65248 14408 65300 14414
rect 65248 14350 65300 14356
rect 65156 7132 65208 7138
rect 65156 7074 65208 7080
rect 65260 5846 65288 14350
rect 65352 11898 65380 22918
rect 65340 11892 65392 11898
rect 65340 11834 65392 11840
rect 65338 11792 65394 11801
rect 65338 11727 65394 11736
rect 65352 7002 65380 11727
rect 65444 9178 65472 24550
rect 65432 9172 65484 9178
rect 65432 9114 65484 9120
rect 65432 9036 65484 9042
rect 65432 8978 65484 8984
rect 65444 7342 65472 8978
rect 65432 7336 65484 7342
rect 65432 7278 65484 7284
rect 65340 6996 65392 7002
rect 65340 6938 65392 6944
rect 65536 6186 65564 28358
rect 65616 26988 65668 26994
rect 65616 26930 65668 26936
rect 65524 6180 65576 6186
rect 65524 6122 65576 6128
rect 65248 5840 65300 5846
rect 65248 5782 65300 5788
rect 65340 5228 65392 5234
rect 65340 5170 65392 5176
rect 65246 5128 65302 5137
rect 65246 5063 65302 5072
rect 65064 4548 65116 4554
rect 65064 4490 65116 4496
rect 65260 4282 65288 5063
rect 65248 4276 65300 4282
rect 65248 4218 65300 4224
rect 65352 4214 65380 5170
rect 65340 4208 65392 4214
rect 64984 4146 65104 4162
rect 65340 4150 65392 4156
rect 64984 4140 65116 4146
rect 64984 4134 65064 4140
rect 64984 3738 65012 4134
rect 65064 4082 65116 4088
rect 65340 3936 65392 3942
rect 65340 3878 65392 3884
rect 64788 3732 64840 3738
rect 64788 3674 64840 3680
rect 64972 3732 65024 3738
rect 64972 3674 65024 3680
rect 64696 2984 64748 2990
rect 64696 2926 64748 2932
rect 64604 2304 64656 2310
rect 64604 2246 64656 2252
rect 64188 2150 64210 2202
rect 64262 2150 64274 2202
rect 64326 2150 64338 2202
rect 64390 2150 64402 2202
rect 64454 2150 64466 2202
rect 64518 2150 64540 2202
rect 64188 1114 64540 2150
rect 64604 1284 64656 1290
rect 64604 1226 64656 1232
rect 64188 1062 64210 1114
rect 64262 1062 64274 1114
rect 64326 1062 64338 1114
rect 64390 1062 64402 1114
rect 64454 1062 64466 1114
rect 64518 1062 64540 1114
rect 64188 1040 64540 1062
rect 64616 1018 64644 1226
rect 64604 1012 64656 1018
rect 64604 954 64656 960
rect 64432 870 64552 898
rect 64432 800 64460 870
rect 54404 734 54616 762
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57058 0 57114 800
rect 57518 0 57574 800
rect 57978 0 58034 800
rect 58438 0 58494 800
rect 58898 0 58954 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60278 0 60334 800
rect 60738 0 60794 800
rect 61198 0 61254 800
rect 61658 0 61714 800
rect 62118 0 62174 800
rect 62578 0 62634 800
rect 63038 0 63094 800
rect 63498 0 63554 800
rect 63958 0 64014 800
rect 64418 0 64474 800
rect 64524 762 64552 870
rect 64708 762 64736 2926
rect 65352 2446 65380 3878
rect 65432 3528 65484 3534
rect 65432 3470 65484 3476
rect 65340 2440 65392 2446
rect 65340 2382 65392 2388
rect 65340 1896 65392 1902
rect 65340 1838 65392 1844
rect 65352 800 65380 1838
rect 65444 1290 65472 3470
rect 65524 2848 65576 2854
rect 65524 2790 65576 2796
rect 65536 2514 65564 2790
rect 65524 2508 65576 2514
rect 65524 2450 65576 2456
rect 65432 1284 65484 1290
rect 65432 1226 65484 1232
rect 65628 1222 65656 26930
rect 65616 1216 65668 1222
rect 65616 1158 65668 1164
rect 64524 734 64736 762
rect 64878 0 64934 800
rect 65338 0 65394 800
rect 65720 134 65748 28426
rect 65812 23866 65840 45902
rect 65984 45620 66036 45626
rect 65984 45562 66036 45568
rect 65892 43648 65944 43654
rect 65892 43590 65944 43596
rect 65904 40934 65932 43590
rect 65892 40928 65944 40934
rect 65892 40870 65944 40876
rect 65892 40724 65944 40730
rect 65892 40666 65944 40672
rect 65904 24410 65932 40666
rect 65996 24410 66024 45562
rect 66088 40730 66116 47058
rect 66076 40724 66128 40730
rect 66076 40666 66128 40672
rect 66076 40588 66128 40594
rect 66076 40530 66128 40536
rect 66088 36174 66116 40530
rect 66180 39642 66208 71606
rect 66352 71596 66404 71602
rect 66352 71538 66404 71544
rect 66260 40928 66312 40934
rect 66260 40870 66312 40876
rect 66168 39636 66220 39642
rect 66168 39578 66220 39584
rect 66272 39522 66300 40870
rect 66364 40730 66392 71538
rect 66628 68672 66680 68678
rect 66628 68614 66680 68620
rect 66536 51536 66588 51542
rect 66536 51478 66588 51484
rect 66444 45280 66496 45286
rect 66444 45222 66496 45228
rect 66352 40724 66404 40730
rect 66352 40666 66404 40672
rect 66352 40180 66404 40186
rect 66352 40122 66404 40128
rect 66180 39494 66300 39522
rect 66076 36168 66128 36174
rect 66076 36110 66128 36116
rect 66180 35986 66208 39494
rect 66088 35958 66208 35986
rect 66088 24818 66116 35958
rect 66364 35894 66392 40122
rect 66180 35866 66392 35894
rect 66180 29850 66208 35866
rect 66168 29844 66220 29850
rect 66168 29786 66220 29792
rect 66352 29640 66404 29646
rect 66352 29582 66404 29588
rect 66260 28008 66312 28014
rect 66260 27950 66312 27956
rect 66076 24812 66128 24818
rect 66076 24754 66128 24760
rect 66168 24744 66220 24750
rect 66168 24686 66220 24692
rect 66076 24608 66128 24614
rect 66076 24550 66128 24556
rect 65892 24404 65944 24410
rect 65892 24346 65944 24352
rect 65984 24404 66036 24410
rect 65984 24346 66036 24352
rect 66088 24206 66116 24550
rect 66076 24200 66128 24206
rect 66076 24142 66128 24148
rect 65892 24064 65944 24070
rect 65892 24006 65944 24012
rect 65800 23860 65852 23866
rect 65800 23802 65852 23808
rect 65904 22094 65932 24006
rect 65812 22066 65932 22094
rect 65812 7410 65840 22066
rect 65892 16788 65944 16794
rect 65892 16730 65944 16736
rect 65800 7404 65852 7410
rect 65800 7346 65852 7352
rect 65904 6458 65932 16730
rect 65984 16652 66036 16658
rect 65984 16594 66036 16600
rect 65996 9042 66024 16594
rect 66088 12753 66116 24142
rect 66180 24070 66208 24686
rect 66168 24064 66220 24070
rect 66168 24006 66220 24012
rect 66168 23792 66220 23798
rect 66168 23734 66220 23740
rect 66074 12744 66130 12753
rect 66074 12679 66130 12688
rect 66076 12640 66128 12646
rect 66076 12582 66128 12588
rect 66088 9217 66116 12582
rect 66074 9208 66130 9217
rect 66074 9143 66130 9152
rect 65984 9036 66036 9042
rect 66180 9024 66208 23734
rect 66272 23254 66300 27950
rect 66260 23248 66312 23254
rect 66260 23190 66312 23196
rect 66260 22568 66312 22574
rect 66260 22510 66312 22516
rect 66272 22409 66300 22510
rect 66258 22400 66314 22409
rect 66258 22335 66314 22344
rect 66260 19168 66312 19174
rect 66260 19110 66312 19116
rect 65984 8978 66036 8984
rect 66088 8996 66208 9024
rect 66088 8922 66116 8996
rect 65996 8894 66116 8922
rect 66166 8936 66222 8945
rect 65996 7274 66024 8894
rect 66166 8871 66222 8880
rect 66076 8832 66128 8838
rect 66076 8774 66128 8780
rect 65984 7268 66036 7274
rect 65984 7210 66036 7216
rect 65892 6452 65944 6458
rect 65892 6394 65944 6400
rect 65892 6180 65944 6186
rect 65892 6122 65944 6128
rect 65800 5840 65852 5846
rect 65800 5782 65852 5788
rect 65812 4049 65840 5782
rect 65904 5642 65932 6122
rect 65892 5636 65944 5642
rect 65892 5578 65944 5584
rect 65984 5364 66036 5370
rect 65984 5306 66036 5312
rect 65798 4040 65854 4049
rect 65798 3975 65854 3984
rect 65892 3460 65944 3466
rect 65892 3402 65944 3408
rect 65904 2650 65932 3402
rect 65892 2644 65944 2650
rect 65892 2586 65944 2592
rect 65800 2508 65852 2514
rect 65800 2450 65852 2456
rect 65812 800 65840 2450
rect 65996 2038 66024 5306
rect 66088 3505 66116 8774
rect 66180 5846 66208 8871
rect 66272 7857 66300 19110
rect 66258 7848 66314 7857
rect 66364 7818 66392 29582
rect 66456 23866 66484 45222
rect 66548 27062 66576 51478
rect 66640 35154 66668 68614
rect 66732 41818 66760 80922
rect 66916 42770 66944 83098
rect 69204 83088 69256 83094
rect 69204 83030 69256 83036
rect 66996 80640 67048 80646
rect 66996 80582 67048 80588
rect 67008 65550 67036 80582
rect 67088 78464 67140 78470
rect 67088 78406 67140 78412
rect 66996 65544 67048 65550
rect 66996 65486 67048 65492
rect 66996 53168 67048 53174
rect 66996 53110 67048 53116
rect 66904 42764 66956 42770
rect 66904 42706 66956 42712
rect 66720 41812 66772 41818
rect 66720 41754 66772 41760
rect 66904 37800 66956 37806
rect 66904 37742 66956 37748
rect 66628 35148 66680 35154
rect 66628 35090 66680 35096
rect 66628 32904 66680 32910
rect 66628 32846 66680 32852
rect 66536 27056 66588 27062
rect 66536 26998 66588 27004
rect 66640 26790 66668 32846
rect 66812 31816 66864 31822
rect 66812 31758 66864 31764
rect 66720 30728 66772 30734
rect 66720 30670 66772 30676
rect 66628 26784 66680 26790
rect 66628 26726 66680 26732
rect 66732 26466 66760 30670
rect 66824 26874 66852 31758
rect 66916 31754 66944 37742
rect 67008 35834 67036 53110
rect 66996 35828 67048 35834
rect 66996 35770 67048 35776
rect 66916 31726 67036 31754
rect 66824 26846 66944 26874
rect 66812 26784 66864 26790
rect 66812 26726 66864 26732
rect 66640 26438 66760 26466
rect 66444 23860 66496 23866
rect 66444 23802 66496 23808
rect 66536 23112 66588 23118
rect 66536 23054 66588 23060
rect 66548 22681 66576 23054
rect 66534 22672 66590 22681
rect 66534 22607 66590 22616
rect 66536 17264 66588 17270
rect 66536 17206 66588 17212
rect 66548 10826 66576 17206
rect 66456 10798 66576 10826
rect 66456 8294 66484 10798
rect 66536 10736 66588 10742
rect 66536 10678 66588 10684
rect 66444 8288 66496 8294
rect 66444 8230 66496 8236
rect 66444 8084 66496 8090
rect 66444 8026 66496 8032
rect 66456 7818 66484 8026
rect 66548 7818 66576 10678
rect 66258 7783 66314 7792
rect 66352 7812 66404 7818
rect 66352 7754 66404 7760
rect 66444 7812 66496 7818
rect 66444 7754 66496 7760
rect 66536 7812 66588 7818
rect 66536 7754 66588 7760
rect 66640 7698 66668 26438
rect 66720 26376 66772 26382
rect 66720 26318 66772 26324
rect 66272 7670 66668 7698
rect 66168 5840 66220 5846
rect 66168 5782 66220 5788
rect 66168 5636 66220 5642
rect 66168 5578 66220 5584
rect 66074 3496 66130 3505
rect 66074 3431 66130 3440
rect 65984 2032 66036 2038
rect 65984 1974 66036 1980
rect 66180 1834 66208 5578
rect 66272 5370 66300 7670
rect 66732 7562 66760 26318
rect 66824 17270 66852 26726
rect 66812 17264 66864 17270
rect 66812 17206 66864 17212
rect 66812 14816 66864 14822
rect 66812 14758 66864 14764
rect 66824 10606 66852 14758
rect 66812 10600 66864 10606
rect 66812 10542 66864 10548
rect 66812 10260 66864 10266
rect 66812 10202 66864 10208
rect 66364 7534 66760 7562
rect 66260 5364 66312 5370
rect 66260 5306 66312 5312
rect 66364 2106 66392 7534
rect 66442 7440 66498 7449
rect 66442 7375 66498 7384
rect 66536 7404 66588 7410
rect 66456 2922 66484 7375
rect 66536 7346 66588 7352
rect 66548 7002 66576 7346
rect 66824 7206 66852 10202
rect 66916 8090 66944 26846
rect 66904 8084 66956 8090
rect 66904 8026 66956 8032
rect 67008 7970 67036 31726
rect 66916 7942 67036 7970
rect 66812 7200 66864 7206
rect 66812 7142 66864 7148
rect 66536 6996 66588 7002
rect 66536 6938 66588 6944
rect 66548 6458 66576 6938
rect 66536 6452 66588 6458
rect 66536 6394 66588 6400
rect 66548 5914 66576 6394
rect 66536 5908 66588 5914
rect 66536 5850 66588 5856
rect 66548 5370 66576 5850
rect 66536 5364 66588 5370
rect 66536 5306 66588 5312
rect 66548 4826 66576 5306
rect 66536 4820 66588 4826
rect 66536 4762 66588 4768
rect 66548 4214 66576 4762
rect 66536 4208 66588 4214
rect 66536 4150 66588 4156
rect 66548 3738 66576 4150
rect 66536 3732 66588 3738
rect 66536 3674 66588 3680
rect 66548 3194 66576 3674
rect 66916 3670 66944 7942
rect 66996 7812 67048 7818
rect 66996 7754 67048 7760
rect 67008 5710 67036 7754
rect 67100 7410 67128 78406
rect 69020 72140 69072 72146
rect 69020 72082 69072 72088
rect 68100 65544 68152 65550
rect 68100 65486 68152 65492
rect 67180 44872 67232 44878
rect 67180 44814 67232 44820
rect 67192 23866 67220 44814
rect 67548 44192 67600 44198
rect 67548 44134 67600 44140
rect 67364 34536 67416 34542
rect 67364 34478 67416 34484
rect 67272 27464 67324 27470
rect 67272 27406 67324 27412
rect 67284 24342 67312 27406
rect 67272 24336 67324 24342
rect 67272 24278 67324 24284
rect 67272 24200 67324 24206
rect 67272 24142 67324 24148
rect 67180 23860 67232 23866
rect 67180 23802 67232 23808
rect 67180 23656 67232 23662
rect 67178 23624 67180 23633
rect 67232 23624 67234 23633
rect 67178 23559 67234 23568
rect 67284 23497 67312 24142
rect 67270 23488 67326 23497
rect 67270 23423 67326 23432
rect 67272 23248 67324 23254
rect 67272 23190 67324 23196
rect 67180 23112 67232 23118
rect 67180 23054 67232 23060
rect 67192 10742 67220 23054
rect 67180 10736 67232 10742
rect 67180 10678 67232 10684
rect 67180 10600 67232 10606
rect 67180 10542 67232 10548
rect 67088 7404 67140 7410
rect 67088 7346 67140 7352
rect 67192 6322 67220 10542
rect 67180 6316 67232 6322
rect 67180 6258 67232 6264
rect 66996 5704 67048 5710
rect 66996 5646 67048 5652
rect 66996 3936 67048 3942
rect 66996 3878 67048 3884
rect 66904 3664 66956 3670
rect 66904 3606 66956 3612
rect 66536 3188 66588 3194
rect 66536 3130 66588 3136
rect 66444 2916 66496 2922
rect 66444 2858 66496 2864
rect 66548 2650 66576 3130
rect 66536 2644 66588 2650
rect 66536 2586 66588 2592
rect 66548 2106 66576 2586
rect 67008 2106 67036 3878
rect 66352 2100 66404 2106
rect 66352 2042 66404 2048
rect 66536 2100 66588 2106
rect 66536 2042 66588 2048
rect 66996 2100 67048 2106
rect 66996 2042 67048 2048
rect 66168 1828 66220 1834
rect 66168 1770 66220 1776
rect 66548 1562 66576 2042
rect 67180 1896 67232 1902
rect 67180 1838 67232 1844
rect 66536 1556 66588 1562
rect 66536 1498 66588 1504
rect 66720 1352 66772 1358
rect 66720 1294 66772 1300
rect 66732 800 66760 1294
rect 67192 800 67220 1838
rect 67284 1494 67312 23190
rect 67376 1766 67404 34478
rect 67456 33992 67508 33998
rect 67456 33934 67508 33940
rect 67468 6866 67496 33934
rect 67560 23322 67588 44134
rect 67916 34604 67968 34610
rect 67916 34546 67968 34552
rect 67640 24336 67692 24342
rect 67640 24278 67692 24284
rect 67548 23316 67600 23322
rect 67548 23258 67600 23264
rect 67652 23202 67680 24278
rect 67732 23656 67784 23662
rect 67732 23598 67784 23604
rect 67560 23174 67680 23202
rect 67456 6860 67508 6866
rect 67456 6802 67508 6808
rect 67560 5642 67588 23174
rect 67640 23112 67692 23118
rect 67640 23054 67692 23060
rect 67652 6225 67680 23054
rect 67744 8090 67772 23598
rect 67824 23588 67876 23594
rect 67824 23530 67876 23536
rect 67836 23118 67864 23530
rect 67824 23112 67876 23118
rect 67824 23054 67876 23060
rect 67824 18964 67876 18970
rect 67824 18906 67876 18912
rect 67732 8084 67784 8090
rect 67732 8026 67784 8032
rect 67836 7970 67864 18906
rect 67744 7942 67864 7970
rect 67928 7954 67956 34546
rect 68008 30184 68060 30190
rect 68008 30126 68060 30132
rect 67916 7948 67968 7954
rect 67638 6216 67694 6225
rect 67638 6151 67694 6160
rect 67548 5636 67600 5642
rect 67548 5578 67600 5584
rect 67744 5574 67772 7942
rect 67916 7890 67968 7896
rect 68020 7834 68048 30126
rect 67836 7806 68048 7834
rect 67836 6361 67864 7806
rect 68112 7698 68140 65486
rect 68560 48136 68612 48142
rect 68560 48078 68612 48084
rect 68376 39432 68428 39438
rect 68376 39374 68428 39380
rect 68192 38344 68244 38350
rect 68192 38286 68244 38292
rect 67928 7670 68140 7698
rect 67822 6352 67878 6361
rect 67822 6287 67878 6296
rect 67732 5568 67784 5574
rect 67732 5510 67784 5516
rect 67928 4146 67956 7670
rect 68204 7562 68232 38286
rect 68284 36168 68336 36174
rect 68284 36110 68336 36116
rect 68020 7534 68232 7562
rect 67916 4140 67968 4146
rect 67916 4082 67968 4088
rect 67928 3738 67956 4082
rect 67916 3732 67968 3738
rect 67916 3674 67968 3680
rect 67548 3596 67600 3602
rect 67548 3538 67600 3544
rect 67364 1760 67416 1766
rect 67364 1702 67416 1708
rect 67272 1488 67324 1494
rect 67272 1430 67324 1436
rect 67560 1290 67588 3538
rect 67640 2984 67692 2990
rect 67640 2926 67692 2932
rect 67652 1358 67680 2926
rect 68020 2038 68048 7534
rect 68100 2848 68152 2854
rect 68100 2790 68152 2796
rect 68112 2446 68140 2790
rect 68100 2440 68152 2446
rect 68100 2382 68152 2388
rect 68008 2032 68060 2038
rect 68008 1974 68060 1980
rect 68296 1562 68324 36110
rect 68388 2514 68416 39374
rect 68468 29776 68520 29782
rect 68468 29718 68520 29724
rect 68480 6662 68508 29718
rect 68468 6656 68520 6662
rect 68468 6598 68520 6604
rect 68572 5681 68600 48078
rect 68652 7948 68704 7954
rect 68652 7890 68704 7896
rect 68558 5672 68614 5681
rect 68558 5607 68614 5616
rect 68664 4865 68692 7890
rect 69032 6186 69060 72082
rect 69112 50380 69164 50386
rect 69112 50322 69164 50328
rect 69020 6180 69072 6186
rect 69020 6122 69072 6128
rect 68650 4856 68706 4865
rect 68650 4791 68706 4800
rect 69124 3398 69152 50322
rect 69216 7546 69244 83030
rect 71836 82236 72188 83206
rect 71836 82180 71864 82236
rect 71920 82180 71944 82236
rect 72000 82180 72024 82236
rect 72080 82180 72104 82236
rect 72160 82180 72188 82236
rect 71836 82170 72188 82180
rect 71836 82118 71858 82170
rect 71910 82156 71922 82170
rect 71974 82156 71986 82170
rect 72038 82156 72050 82170
rect 72102 82156 72114 82170
rect 71920 82118 71922 82156
rect 72102 82118 72104 82156
rect 72166 82118 72188 82170
rect 71836 82100 71864 82118
rect 71920 82100 71944 82118
rect 72000 82100 72024 82118
rect 72080 82100 72104 82118
rect 72160 82100 72188 82118
rect 71836 82076 72188 82100
rect 71836 82020 71864 82076
rect 71920 82020 71944 82076
rect 72000 82020 72024 82076
rect 72080 82020 72104 82076
rect 72160 82020 72188 82076
rect 71836 81996 72188 82020
rect 71836 81940 71864 81996
rect 71920 81940 71944 81996
rect 72000 81940 72024 81996
rect 72080 81940 72104 81996
rect 72160 81940 72188 81996
rect 71836 81082 72188 81940
rect 71836 81030 71858 81082
rect 71910 81030 71922 81082
rect 71974 81030 71986 81082
rect 72038 81030 72050 81082
rect 72102 81030 72114 81082
rect 72166 81030 72188 81082
rect 71836 79994 72188 81030
rect 71836 79942 71858 79994
rect 71910 79942 71922 79994
rect 71974 79942 71986 79994
rect 72038 79942 72050 79994
rect 72102 79942 72114 79994
rect 72166 79942 72188 79994
rect 71836 78906 72188 79942
rect 71836 78854 71858 78906
rect 71910 78854 71922 78906
rect 71974 78854 71986 78906
rect 72038 78854 72050 78906
rect 72102 78854 72114 78906
rect 72166 78854 72188 78906
rect 71836 77818 72188 78854
rect 71836 77766 71858 77818
rect 71910 77766 71922 77818
rect 71974 77766 71986 77818
rect 72038 77766 72050 77818
rect 72102 77766 72114 77818
rect 72166 77766 72188 77818
rect 71836 76730 72188 77766
rect 71836 76678 71858 76730
rect 71910 76678 71922 76730
rect 71974 76678 71986 76730
rect 72038 76678 72050 76730
rect 72102 76678 72114 76730
rect 72166 76678 72188 76730
rect 71836 75642 72188 76678
rect 71836 75590 71858 75642
rect 71910 75590 71922 75642
rect 71974 75590 71986 75642
rect 72038 75590 72050 75642
rect 72102 75590 72114 75642
rect 72166 75590 72188 75642
rect 71836 74554 72188 75590
rect 71836 74502 71858 74554
rect 71910 74502 71922 74554
rect 71974 74502 71986 74554
rect 72038 74502 72050 74554
rect 72102 74502 72114 74554
rect 72166 74502 72188 74554
rect 71836 73466 72188 74502
rect 71836 73414 71858 73466
rect 71910 73414 71922 73466
rect 71974 73414 71986 73466
rect 72038 73414 72050 73466
rect 72102 73414 72114 73466
rect 72166 73414 72188 73466
rect 71836 72378 72188 73414
rect 71836 72326 71858 72378
rect 71910 72326 71922 72378
rect 71974 72326 71986 72378
rect 72038 72326 72050 72378
rect 72102 72326 72114 72378
rect 72166 72326 72188 72378
rect 71836 72236 72188 72326
rect 71836 72180 71864 72236
rect 71920 72180 71944 72236
rect 72000 72180 72024 72236
rect 72080 72180 72104 72236
rect 72160 72180 72188 72236
rect 71836 72156 72188 72180
rect 71836 72100 71864 72156
rect 71920 72100 71944 72156
rect 72000 72100 72024 72156
rect 72080 72100 72104 72156
rect 72160 72100 72188 72156
rect 71836 72076 72188 72100
rect 71836 72020 71864 72076
rect 71920 72020 71944 72076
rect 72000 72020 72024 72076
rect 72080 72020 72104 72076
rect 72160 72020 72188 72076
rect 71836 71996 72188 72020
rect 71836 71940 71864 71996
rect 71920 71940 71944 71996
rect 72000 71940 72024 71996
rect 72080 71940 72104 71996
rect 72160 71940 72188 71996
rect 71836 71290 72188 71940
rect 71836 71238 71858 71290
rect 71910 71238 71922 71290
rect 71974 71238 71986 71290
rect 72038 71238 72050 71290
rect 72102 71238 72114 71290
rect 72166 71238 72188 71290
rect 71836 70202 72188 71238
rect 71836 70150 71858 70202
rect 71910 70150 71922 70202
rect 71974 70150 71986 70202
rect 72038 70150 72050 70202
rect 72102 70150 72114 70202
rect 72166 70150 72188 70202
rect 71836 69114 72188 70150
rect 71836 69062 71858 69114
rect 71910 69062 71922 69114
rect 71974 69062 71986 69114
rect 72038 69062 72050 69114
rect 72102 69062 72114 69114
rect 72166 69062 72188 69114
rect 71836 68026 72188 69062
rect 71836 67974 71858 68026
rect 71910 67974 71922 68026
rect 71974 67974 71986 68026
rect 72038 67974 72050 68026
rect 72102 67974 72114 68026
rect 72166 67974 72188 68026
rect 71836 66938 72188 67974
rect 71836 66886 71858 66938
rect 71910 66886 71922 66938
rect 71974 66886 71986 66938
rect 72038 66886 72050 66938
rect 72102 66886 72114 66938
rect 72166 66886 72188 66938
rect 71836 65850 72188 66886
rect 71836 65798 71858 65850
rect 71910 65798 71922 65850
rect 71974 65798 71986 65850
rect 72038 65798 72050 65850
rect 72102 65798 72114 65850
rect 72166 65798 72188 65850
rect 71836 64762 72188 65798
rect 71836 64710 71858 64762
rect 71910 64710 71922 64762
rect 71974 64710 71986 64762
rect 72038 64710 72050 64762
rect 72102 64710 72114 64762
rect 72166 64710 72188 64762
rect 71836 63674 72188 64710
rect 71836 63622 71858 63674
rect 71910 63622 71922 63674
rect 71974 63622 71986 63674
rect 72038 63622 72050 63674
rect 72102 63622 72114 63674
rect 72166 63622 72188 63674
rect 71836 62586 72188 63622
rect 71836 62534 71858 62586
rect 71910 62534 71922 62586
rect 71974 62534 71986 62586
rect 72038 62534 72050 62586
rect 72102 62534 72114 62586
rect 72166 62534 72188 62586
rect 71836 62236 72188 62534
rect 71836 62180 71864 62236
rect 71920 62180 71944 62236
rect 72000 62180 72024 62236
rect 72080 62180 72104 62236
rect 72160 62180 72188 62236
rect 71836 62156 72188 62180
rect 71836 62100 71864 62156
rect 71920 62100 71944 62156
rect 72000 62100 72024 62156
rect 72080 62100 72104 62156
rect 72160 62100 72188 62156
rect 71836 62076 72188 62100
rect 71836 62020 71864 62076
rect 71920 62020 71944 62076
rect 72000 62020 72024 62076
rect 72080 62020 72104 62076
rect 72160 62020 72188 62076
rect 71836 61996 72188 62020
rect 71836 61940 71864 61996
rect 71920 61940 71944 61996
rect 72000 61940 72024 61996
rect 72080 61940 72104 61996
rect 72160 61940 72188 61996
rect 71836 61498 72188 61940
rect 71836 61446 71858 61498
rect 71910 61446 71922 61498
rect 71974 61446 71986 61498
rect 72038 61446 72050 61498
rect 72102 61446 72114 61498
rect 72166 61446 72188 61498
rect 71836 60410 72188 61446
rect 71836 60358 71858 60410
rect 71910 60358 71922 60410
rect 71974 60358 71986 60410
rect 72038 60358 72050 60410
rect 72102 60358 72114 60410
rect 72166 60358 72188 60410
rect 71836 59322 72188 60358
rect 71836 59270 71858 59322
rect 71910 59270 71922 59322
rect 71974 59270 71986 59322
rect 72038 59270 72050 59322
rect 72102 59270 72114 59322
rect 72166 59270 72188 59322
rect 71836 58234 72188 59270
rect 71836 58182 71858 58234
rect 71910 58182 71922 58234
rect 71974 58182 71986 58234
rect 72038 58182 72050 58234
rect 72102 58182 72114 58234
rect 72166 58182 72188 58234
rect 71836 57146 72188 58182
rect 71836 57094 71858 57146
rect 71910 57094 71922 57146
rect 71974 57094 71986 57146
rect 72038 57094 72050 57146
rect 72102 57094 72114 57146
rect 72166 57094 72188 57146
rect 71836 56058 72188 57094
rect 71836 56006 71858 56058
rect 71910 56006 71922 56058
rect 71974 56006 71986 56058
rect 72038 56006 72050 56058
rect 72102 56006 72114 56058
rect 72166 56006 72188 56058
rect 71836 54970 72188 56006
rect 71836 54918 71858 54970
rect 71910 54918 71922 54970
rect 71974 54918 71986 54970
rect 72038 54918 72050 54970
rect 72102 54918 72114 54970
rect 72166 54918 72188 54970
rect 71836 53882 72188 54918
rect 71836 53830 71858 53882
rect 71910 53830 71922 53882
rect 71974 53830 71986 53882
rect 72038 53830 72050 53882
rect 72102 53830 72114 53882
rect 72166 53830 72188 53882
rect 71836 52794 72188 53830
rect 71836 52742 71858 52794
rect 71910 52742 71922 52794
rect 71974 52742 71986 52794
rect 72038 52742 72050 52794
rect 72102 52742 72114 52794
rect 72166 52742 72188 52794
rect 69296 52624 69348 52630
rect 69296 52566 69348 52572
rect 69204 7540 69256 7546
rect 69204 7482 69256 7488
rect 69216 7002 69244 7482
rect 69204 6996 69256 7002
rect 69204 6938 69256 6944
rect 69216 6458 69244 6938
rect 69308 6798 69336 52566
rect 71836 52236 72188 52742
rect 71836 52180 71864 52236
rect 71920 52180 71944 52236
rect 72000 52180 72024 52236
rect 72080 52180 72104 52236
rect 72160 52180 72188 52236
rect 71836 52156 72188 52180
rect 71836 52100 71864 52156
rect 71920 52100 71944 52156
rect 72000 52100 72024 52156
rect 72080 52100 72104 52156
rect 72160 52100 72188 52156
rect 71836 52076 72188 52100
rect 71836 52020 71864 52076
rect 71920 52020 71944 52076
rect 72000 52020 72024 52076
rect 72080 52020 72104 52076
rect 72160 52020 72188 52076
rect 71836 51996 72188 52020
rect 71836 51940 71864 51996
rect 71920 51940 71944 51996
rect 72000 51940 72024 51996
rect 72080 51940 72104 51996
rect 72160 51940 72188 51996
rect 71836 51706 72188 51940
rect 71836 51654 71858 51706
rect 71910 51654 71922 51706
rect 71974 51654 71986 51706
rect 72038 51654 72050 51706
rect 72102 51654 72114 51706
rect 72166 51654 72188 51706
rect 71836 50618 72188 51654
rect 71836 50566 71858 50618
rect 71910 50566 71922 50618
rect 71974 50566 71986 50618
rect 72038 50566 72050 50618
rect 72102 50566 72114 50618
rect 72166 50566 72188 50618
rect 71836 49530 72188 50566
rect 71836 49478 71858 49530
rect 71910 49478 71922 49530
rect 71974 49478 71986 49530
rect 72038 49478 72050 49530
rect 72102 49478 72114 49530
rect 72166 49478 72188 49530
rect 71836 48442 72188 49478
rect 71836 48390 71858 48442
rect 71910 48390 71922 48442
rect 71974 48390 71986 48442
rect 72038 48390 72050 48442
rect 72102 48390 72114 48442
rect 72166 48390 72188 48442
rect 71836 47354 72188 48390
rect 71836 47302 71858 47354
rect 71910 47302 71922 47354
rect 71974 47302 71986 47354
rect 72038 47302 72050 47354
rect 72102 47302 72114 47354
rect 72166 47302 72188 47354
rect 71836 46266 72188 47302
rect 71836 46214 71858 46266
rect 71910 46214 71922 46266
rect 71974 46214 71986 46266
rect 72038 46214 72050 46266
rect 72102 46214 72114 46266
rect 72166 46214 72188 46266
rect 71836 45178 72188 46214
rect 71836 45126 71858 45178
rect 71910 45126 71922 45178
rect 71974 45126 71986 45178
rect 72038 45126 72050 45178
rect 72102 45126 72114 45178
rect 72166 45126 72188 45178
rect 71836 44090 72188 45126
rect 71836 44038 71858 44090
rect 71910 44038 71922 44090
rect 71974 44038 71986 44090
rect 72038 44038 72050 44090
rect 72102 44038 72114 44090
rect 72166 44038 72188 44090
rect 69388 43308 69440 43314
rect 69388 43250 69440 43256
rect 69296 6792 69348 6798
rect 69296 6734 69348 6740
rect 69204 6452 69256 6458
rect 69204 6394 69256 6400
rect 69216 5914 69244 6394
rect 69400 6390 69428 43250
rect 71836 43002 72188 44038
rect 71836 42950 71858 43002
rect 71910 42950 71922 43002
rect 71974 42950 71986 43002
rect 72038 42950 72050 43002
rect 72102 42950 72114 43002
rect 72166 42950 72188 43002
rect 69664 42696 69716 42702
rect 69664 42638 69716 42644
rect 69480 40656 69532 40662
rect 69480 40598 69532 40604
rect 69388 6384 69440 6390
rect 69388 6326 69440 6332
rect 69204 5908 69256 5914
rect 69204 5850 69256 5856
rect 69216 5370 69244 5850
rect 69492 5817 69520 40598
rect 69572 32428 69624 32434
rect 69572 32370 69624 32376
rect 69584 6118 69612 32370
rect 69572 6112 69624 6118
rect 69572 6054 69624 6060
rect 69478 5808 69534 5817
rect 69478 5743 69534 5752
rect 69204 5364 69256 5370
rect 69204 5306 69256 5312
rect 69216 4826 69244 5306
rect 69204 4820 69256 4826
rect 69204 4762 69256 4768
rect 69216 4214 69244 4762
rect 69204 4208 69256 4214
rect 69204 4150 69256 4156
rect 69216 3738 69244 4150
rect 69388 3936 69440 3942
rect 69388 3878 69440 3884
rect 69204 3732 69256 3738
rect 69204 3674 69256 3680
rect 69112 3392 69164 3398
rect 69112 3334 69164 3340
rect 69216 3194 69244 3674
rect 69204 3188 69256 3194
rect 69204 3130 69256 3136
rect 68560 2984 68612 2990
rect 68560 2926 68612 2932
rect 68376 2508 68428 2514
rect 68376 2450 68428 2456
rect 68284 1556 68336 1562
rect 68284 1498 68336 1504
rect 67640 1352 67692 1358
rect 67640 1294 67692 1300
rect 68100 1352 68152 1358
rect 68100 1294 68152 1300
rect 67548 1284 67600 1290
rect 67548 1226 67600 1232
rect 68112 800 68140 1294
rect 68572 800 68600 2926
rect 69216 2650 69244 3130
rect 69400 3058 69428 3878
rect 69388 3052 69440 3058
rect 69388 2994 69440 3000
rect 69204 2644 69256 2650
rect 69204 2586 69256 2592
rect 69216 2038 69244 2586
rect 69480 2440 69532 2446
rect 69480 2382 69532 2388
rect 69204 2032 69256 2038
rect 69204 1974 69256 1980
rect 69216 1562 69244 1974
rect 69388 1828 69440 1834
rect 69388 1770 69440 1776
rect 69204 1556 69256 1562
rect 69204 1498 69256 1504
rect 69400 1000 69428 1770
rect 69492 1562 69520 2382
rect 69676 2378 69704 42638
rect 71836 42236 72188 42950
rect 71836 42180 71864 42236
rect 71920 42180 71944 42236
rect 72000 42180 72024 42236
rect 72080 42180 72104 42236
rect 72160 42180 72188 42236
rect 71836 42156 72188 42180
rect 71836 42100 71864 42156
rect 71920 42100 71944 42156
rect 72000 42100 72024 42156
rect 72080 42100 72104 42156
rect 72160 42100 72188 42156
rect 71836 42076 72188 42100
rect 71836 42020 71864 42076
rect 71920 42020 71944 42076
rect 72000 42020 72024 42076
rect 72080 42020 72104 42076
rect 72160 42020 72188 42076
rect 71836 41996 72188 42020
rect 71836 41940 71864 41996
rect 71920 41940 71944 41996
rect 72000 41940 72024 41996
rect 72080 41940 72104 41996
rect 72160 41940 72188 41996
rect 71836 41914 72188 41940
rect 71836 41862 71858 41914
rect 71910 41862 71922 41914
rect 71974 41862 71986 41914
rect 72038 41862 72050 41914
rect 72102 41862 72114 41914
rect 72166 41862 72188 41914
rect 69848 41608 69900 41614
rect 69848 41550 69900 41556
rect 69860 2514 69888 41550
rect 71836 40826 72188 41862
rect 71836 40774 71858 40826
rect 71910 40774 71922 40826
rect 71974 40774 71986 40826
rect 72038 40774 72050 40826
rect 72102 40774 72114 40826
rect 72166 40774 72188 40826
rect 70032 40520 70084 40526
rect 70032 40462 70084 40468
rect 69940 25696 69992 25702
rect 69940 25638 69992 25644
rect 69952 3641 69980 25638
rect 69938 3632 69994 3641
rect 69938 3567 69994 3576
rect 69848 2508 69900 2514
rect 69848 2450 69900 2456
rect 69664 2372 69716 2378
rect 69664 2314 69716 2320
rect 70044 2038 70072 40462
rect 71836 39738 72188 40774
rect 71836 39686 71858 39738
rect 71910 39686 71922 39738
rect 71974 39686 71986 39738
rect 72038 39686 72050 39738
rect 72102 39686 72114 39738
rect 72166 39686 72188 39738
rect 71836 38650 72188 39686
rect 71836 38598 71858 38650
rect 71910 38598 71922 38650
rect 71974 38598 71986 38650
rect 72038 38598 72050 38650
rect 72102 38598 72114 38650
rect 72166 38598 72188 38650
rect 71836 37562 72188 38598
rect 71836 37510 71858 37562
rect 71910 37510 71922 37562
rect 71974 37510 71986 37562
rect 72038 37510 72050 37562
rect 72102 37510 72114 37562
rect 72166 37510 72188 37562
rect 71836 36474 72188 37510
rect 71836 36422 71858 36474
rect 71910 36422 71922 36474
rect 71974 36422 71986 36474
rect 72038 36422 72050 36474
rect 72102 36422 72114 36474
rect 72166 36422 72188 36474
rect 71836 35386 72188 36422
rect 71836 35334 71858 35386
rect 71910 35334 71922 35386
rect 71974 35334 71986 35386
rect 72038 35334 72050 35386
rect 72102 35334 72114 35386
rect 72166 35334 72188 35386
rect 71836 34298 72188 35334
rect 71836 34246 71858 34298
rect 71910 34246 71922 34298
rect 71974 34246 71986 34298
rect 72038 34246 72050 34298
rect 72102 34246 72114 34298
rect 72166 34246 72188 34298
rect 71836 33210 72188 34246
rect 71836 33158 71858 33210
rect 71910 33158 71922 33210
rect 71974 33158 71986 33210
rect 72038 33158 72050 33210
rect 72102 33158 72114 33210
rect 72166 33158 72188 33210
rect 71836 32236 72188 33158
rect 71836 32180 71864 32236
rect 71920 32180 71944 32236
rect 72000 32180 72024 32236
rect 72080 32180 72104 32236
rect 72160 32180 72188 32236
rect 71836 32156 72188 32180
rect 71836 32122 71864 32156
rect 71920 32122 71944 32156
rect 72000 32122 72024 32156
rect 72080 32122 72104 32156
rect 72160 32122 72188 32156
rect 71836 32070 71858 32122
rect 71920 32100 71922 32122
rect 72102 32100 72104 32122
rect 71910 32076 71922 32100
rect 71974 32076 71986 32100
rect 72038 32076 72050 32100
rect 72102 32076 72114 32100
rect 71920 32070 71922 32076
rect 72102 32070 72104 32076
rect 72166 32070 72188 32122
rect 71836 32020 71864 32070
rect 71920 32020 71944 32070
rect 72000 32020 72024 32070
rect 72080 32020 72104 32070
rect 72160 32020 72188 32070
rect 71836 31996 72188 32020
rect 71836 31940 71864 31996
rect 71920 31940 71944 31996
rect 72000 31940 72024 31996
rect 72080 31940 72104 31996
rect 72160 31940 72188 31996
rect 71836 31034 72188 31940
rect 71836 30982 71858 31034
rect 71910 30982 71922 31034
rect 71974 30982 71986 31034
rect 72038 30982 72050 31034
rect 72102 30982 72114 31034
rect 72166 30982 72188 31034
rect 71836 29946 72188 30982
rect 71836 29894 71858 29946
rect 71910 29894 71922 29946
rect 71974 29894 71986 29946
rect 72038 29894 72050 29946
rect 72102 29894 72114 29946
rect 72166 29894 72188 29946
rect 71836 28858 72188 29894
rect 71836 28806 71858 28858
rect 71910 28806 71922 28858
rect 71974 28806 71986 28858
rect 72038 28806 72050 28858
rect 72102 28806 72114 28858
rect 72166 28806 72188 28858
rect 70124 27872 70176 27878
rect 70124 27814 70176 27820
rect 70136 4486 70164 27814
rect 71836 27770 72188 28806
rect 71836 27718 71858 27770
rect 71910 27718 71922 27770
rect 71974 27718 71986 27770
rect 72038 27718 72050 27770
rect 72102 27718 72114 27770
rect 72166 27718 72188 27770
rect 71836 26682 72188 27718
rect 71836 26630 71858 26682
rect 71910 26630 71922 26682
rect 71974 26630 71986 26682
rect 72038 26630 72050 26682
rect 72102 26630 72114 26682
rect 72166 26630 72188 26682
rect 71836 25594 72188 26630
rect 71836 25542 71858 25594
rect 71910 25542 71922 25594
rect 71974 25542 71986 25594
rect 72038 25542 72050 25594
rect 72102 25542 72114 25594
rect 72166 25542 72188 25594
rect 71836 24506 72188 25542
rect 71836 24454 71858 24506
rect 71910 24454 71922 24506
rect 71974 24454 71986 24506
rect 72038 24454 72050 24506
rect 72102 24454 72114 24506
rect 72166 24454 72188 24506
rect 71836 23418 72188 24454
rect 71836 23366 71858 23418
rect 71910 23366 71922 23418
rect 71974 23366 71986 23418
rect 72038 23366 72050 23418
rect 72102 23366 72114 23418
rect 72166 23366 72188 23418
rect 71836 22330 72188 23366
rect 71836 22278 71858 22330
rect 71910 22278 71922 22330
rect 71974 22278 71986 22330
rect 72038 22278 72050 22330
rect 72102 22278 72114 22330
rect 72166 22278 72188 22330
rect 71836 22236 72188 22278
rect 71836 22180 71864 22236
rect 71920 22180 71944 22236
rect 72000 22180 72024 22236
rect 72080 22180 72104 22236
rect 72160 22180 72188 22236
rect 71836 22156 72188 22180
rect 71836 22100 71864 22156
rect 71920 22100 71944 22156
rect 72000 22100 72024 22156
rect 72080 22100 72104 22156
rect 72160 22100 72188 22156
rect 71836 22076 72188 22100
rect 71836 22020 71864 22076
rect 71920 22020 71944 22076
rect 72000 22020 72024 22076
rect 72080 22020 72104 22076
rect 72160 22020 72188 22076
rect 71836 21996 72188 22020
rect 71836 21940 71864 21996
rect 71920 21940 71944 21996
rect 72000 21940 72024 21996
rect 72080 21940 72104 21996
rect 72160 21940 72188 21996
rect 70216 21412 70268 21418
rect 70216 21354 70268 21360
rect 70228 5778 70256 21354
rect 71836 21242 72188 21940
rect 71836 21190 71858 21242
rect 71910 21190 71922 21242
rect 71974 21190 71986 21242
rect 72038 21190 72050 21242
rect 72102 21190 72114 21242
rect 72166 21190 72188 21242
rect 71836 20154 72188 21190
rect 71836 20102 71858 20154
rect 71910 20102 71922 20154
rect 71974 20102 71986 20154
rect 72038 20102 72050 20154
rect 72102 20102 72114 20154
rect 72166 20102 72188 20154
rect 71836 19066 72188 20102
rect 71836 19014 71858 19066
rect 71910 19014 71922 19066
rect 71974 19014 71986 19066
rect 72038 19014 72050 19066
rect 72102 19014 72114 19066
rect 72166 19014 72188 19066
rect 71836 17978 72188 19014
rect 71836 17926 71858 17978
rect 71910 17926 71922 17978
rect 71974 17926 71986 17978
rect 72038 17926 72050 17978
rect 72102 17926 72114 17978
rect 72166 17926 72188 17978
rect 71836 16890 72188 17926
rect 71836 16838 71858 16890
rect 71910 16838 71922 16890
rect 71974 16838 71986 16890
rect 72038 16838 72050 16890
rect 72102 16838 72114 16890
rect 72166 16838 72188 16890
rect 71836 15802 72188 16838
rect 71836 15750 71858 15802
rect 71910 15750 71922 15802
rect 71974 15750 71986 15802
rect 72038 15750 72050 15802
rect 72102 15750 72114 15802
rect 72166 15750 72188 15802
rect 71836 14714 72188 15750
rect 71836 14662 71858 14714
rect 71910 14662 71922 14714
rect 71974 14662 71986 14714
rect 72038 14662 72050 14714
rect 72102 14662 72114 14714
rect 72166 14662 72188 14714
rect 71836 13626 72188 14662
rect 71836 13574 71858 13626
rect 71910 13574 71922 13626
rect 71974 13574 71986 13626
rect 72038 13574 72050 13626
rect 72102 13574 72114 13626
rect 72166 13574 72188 13626
rect 71836 12538 72188 13574
rect 71836 12486 71858 12538
rect 71910 12486 71922 12538
rect 71974 12486 71986 12538
rect 72038 12486 72050 12538
rect 72102 12486 72114 12538
rect 72166 12486 72188 12538
rect 71836 12236 72188 12486
rect 71836 12180 71864 12236
rect 71920 12180 71944 12236
rect 72000 12180 72024 12236
rect 72080 12180 72104 12236
rect 72160 12180 72188 12236
rect 71836 12156 72188 12180
rect 71836 12100 71864 12156
rect 71920 12100 71944 12156
rect 72000 12100 72024 12156
rect 72080 12100 72104 12156
rect 72160 12100 72188 12156
rect 71836 12076 72188 12100
rect 71836 12020 71864 12076
rect 71920 12020 71944 12076
rect 72000 12020 72024 12076
rect 72080 12020 72104 12076
rect 72160 12020 72188 12076
rect 71836 11996 72188 12020
rect 71836 11940 71864 11996
rect 71920 11940 71944 11996
rect 72000 11940 72024 11996
rect 72080 11940 72104 11996
rect 72160 11940 72188 11996
rect 71836 11450 72188 11940
rect 71836 11398 71858 11450
rect 71910 11398 71922 11450
rect 71974 11398 71986 11450
rect 72038 11398 72050 11450
rect 72102 11398 72114 11450
rect 72166 11398 72188 11450
rect 71836 10362 72188 11398
rect 71836 10310 71858 10362
rect 71910 10310 71922 10362
rect 71974 10310 71986 10362
rect 72038 10310 72050 10362
rect 72102 10310 72114 10362
rect 72166 10310 72188 10362
rect 71836 9274 72188 10310
rect 71836 9222 71858 9274
rect 71910 9222 71922 9274
rect 71974 9222 71986 9274
rect 72038 9222 72050 9274
rect 72102 9222 72114 9274
rect 72166 9222 72188 9274
rect 71836 8186 72188 9222
rect 71836 8134 71858 8186
rect 71910 8134 71922 8186
rect 71974 8134 71986 8186
rect 72038 8134 72050 8186
rect 72102 8134 72114 8186
rect 72166 8134 72188 8186
rect 71836 7098 72188 8134
rect 71836 7046 71858 7098
rect 71910 7046 71922 7098
rect 71974 7046 71986 7098
rect 72038 7046 72050 7098
rect 72102 7046 72114 7098
rect 72166 7046 72188 7098
rect 71836 6010 72188 7046
rect 71836 5958 71858 6010
rect 71910 5958 71922 6010
rect 71974 5958 71986 6010
rect 72038 5958 72050 6010
rect 72102 5958 72114 6010
rect 72166 5958 72188 6010
rect 70216 5772 70268 5778
rect 70216 5714 70268 5720
rect 71836 4922 72188 5958
rect 71836 4870 71858 4922
rect 71910 4870 71922 4922
rect 71974 4870 71986 4922
rect 72038 4870 72050 4922
rect 72102 4870 72114 4922
rect 72166 4870 72188 4922
rect 70124 4480 70176 4486
rect 70124 4422 70176 4428
rect 70584 4004 70636 4010
rect 70584 3946 70636 3952
rect 70032 2032 70084 2038
rect 70032 1974 70084 1980
rect 69480 1556 69532 1562
rect 69480 1498 69532 1504
rect 69940 1420 69992 1426
rect 69940 1362 69992 1368
rect 69400 972 69520 1000
rect 69492 800 69520 972
rect 69952 800 69980 1362
rect 70596 1358 70624 3946
rect 71412 3936 71464 3942
rect 71412 3878 71464 3884
rect 70676 2440 70728 2446
rect 70676 2382 70728 2388
rect 70688 2106 70716 2382
rect 70860 2304 70912 2310
rect 70860 2246 70912 2252
rect 70676 2100 70728 2106
rect 70676 2042 70728 2048
rect 70872 1970 70900 2246
rect 71424 1970 71452 3878
rect 71836 3834 72188 4870
rect 71836 3782 71858 3834
rect 71910 3782 71922 3834
rect 71974 3782 71986 3834
rect 72038 3782 72050 3834
rect 72102 3782 72114 3834
rect 72166 3782 72188 3834
rect 71836 2746 72188 3782
rect 71836 2694 71858 2746
rect 71910 2694 71922 2746
rect 71974 2694 71986 2746
rect 72038 2694 72050 2746
rect 72102 2694 72114 2746
rect 72166 2694 72188 2746
rect 71836 2236 72188 2694
rect 74188 85978 74540 86000
rect 74188 85926 74210 85978
rect 74262 85926 74274 85978
rect 74326 85926 74338 85978
rect 74390 85926 74402 85978
rect 74454 85926 74466 85978
rect 74518 85926 74540 85978
rect 74188 84890 74540 85926
rect 74188 84838 74210 84890
rect 74262 84838 74274 84890
rect 74326 84838 74338 84890
rect 74390 84838 74402 84890
rect 74454 84838 74466 84890
rect 74518 84838 74540 84890
rect 74188 84588 74540 84838
rect 74188 84532 74216 84588
rect 74272 84532 74296 84588
rect 74352 84532 74376 84588
rect 74432 84532 74456 84588
rect 74512 84532 74540 84588
rect 74188 84508 74540 84532
rect 74188 84452 74216 84508
rect 74272 84452 74296 84508
rect 74352 84452 74376 84508
rect 74432 84452 74456 84508
rect 74512 84452 74540 84508
rect 74188 84428 74540 84452
rect 74188 84372 74216 84428
rect 74272 84372 74296 84428
rect 74352 84372 74376 84428
rect 74432 84372 74456 84428
rect 74512 84372 74540 84428
rect 74188 84348 74540 84372
rect 74188 84292 74216 84348
rect 74272 84292 74296 84348
rect 74352 84292 74376 84348
rect 74432 84292 74456 84348
rect 74512 84292 74540 84348
rect 74188 83802 74540 84292
rect 74188 83750 74210 83802
rect 74262 83750 74274 83802
rect 74326 83750 74338 83802
rect 74390 83750 74402 83802
rect 74454 83750 74466 83802
rect 74518 83750 74540 83802
rect 74188 82714 74540 83750
rect 74188 82662 74210 82714
rect 74262 82662 74274 82714
rect 74326 82662 74338 82714
rect 74390 82662 74402 82714
rect 74454 82662 74466 82714
rect 74518 82662 74540 82714
rect 74188 81626 74540 82662
rect 74188 81574 74210 81626
rect 74262 81574 74274 81626
rect 74326 81574 74338 81626
rect 74390 81574 74402 81626
rect 74454 81574 74466 81626
rect 74518 81574 74540 81626
rect 74188 80538 74540 81574
rect 74188 80486 74210 80538
rect 74262 80486 74274 80538
rect 74326 80486 74338 80538
rect 74390 80486 74402 80538
rect 74454 80486 74466 80538
rect 74518 80486 74540 80538
rect 74188 79450 74540 80486
rect 74188 79398 74210 79450
rect 74262 79398 74274 79450
rect 74326 79398 74338 79450
rect 74390 79398 74402 79450
rect 74454 79398 74466 79450
rect 74518 79398 74540 79450
rect 74188 78362 74540 79398
rect 74188 78310 74210 78362
rect 74262 78310 74274 78362
rect 74326 78310 74338 78362
rect 74390 78310 74402 78362
rect 74454 78310 74466 78362
rect 74518 78310 74540 78362
rect 74188 77274 74540 78310
rect 74188 77222 74210 77274
rect 74262 77222 74274 77274
rect 74326 77222 74338 77274
rect 74390 77222 74402 77274
rect 74454 77222 74466 77274
rect 74518 77222 74540 77274
rect 74188 76186 74540 77222
rect 74188 76134 74210 76186
rect 74262 76134 74274 76186
rect 74326 76134 74338 76186
rect 74390 76134 74402 76186
rect 74454 76134 74466 76186
rect 74518 76134 74540 76186
rect 74188 75098 74540 76134
rect 74188 75046 74210 75098
rect 74262 75046 74274 75098
rect 74326 75046 74338 75098
rect 74390 75046 74402 75098
rect 74454 75046 74466 75098
rect 74518 75046 74540 75098
rect 74188 74588 74540 75046
rect 74188 74532 74216 74588
rect 74272 74532 74296 74588
rect 74352 74532 74376 74588
rect 74432 74532 74456 74588
rect 74512 74532 74540 74588
rect 74188 74508 74540 74532
rect 74188 74452 74216 74508
rect 74272 74452 74296 74508
rect 74352 74452 74376 74508
rect 74432 74452 74456 74508
rect 74512 74452 74540 74508
rect 74188 74428 74540 74452
rect 74188 74372 74216 74428
rect 74272 74372 74296 74428
rect 74352 74372 74376 74428
rect 74432 74372 74456 74428
rect 74512 74372 74540 74428
rect 74188 74348 74540 74372
rect 74188 74292 74216 74348
rect 74272 74292 74296 74348
rect 74352 74292 74376 74348
rect 74432 74292 74456 74348
rect 74512 74292 74540 74348
rect 74188 74010 74540 74292
rect 74188 73958 74210 74010
rect 74262 73958 74274 74010
rect 74326 73958 74338 74010
rect 74390 73958 74402 74010
rect 74454 73958 74466 74010
rect 74518 73958 74540 74010
rect 74188 72922 74540 73958
rect 74188 72870 74210 72922
rect 74262 72870 74274 72922
rect 74326 72870 74338 72922
rect 74390 72870 74402 72922
rect 74454 72870 74466 72922
rect 74518 72870 74540 72922
rect 74188 71834 74540 72870
rect 74188 71782 74210 71834
rect 74262 71782 74274 71834
rect 74326 71782 74338 71834
rect 74390 71782 74402 71834
rect 74454 71782 74466 71834
rect 74518 71782 74540 71834
rect 74188 70746 74540 71782
rect 74188 70694 74210 70746
rect 74262 70694 74274 70746
rect 74326 70694 74338 70746
rect 74390 70694 74402 70746
rect 74454 70694 74466 70746
rect 74518 70694 74540 70746
rect 74188 69658 74540 70694
rect 74188 69606 74210 69658
rect 74262 69606 74274 69658
rect 74326 69606 74338 69658
rect 74390 69606 74402 69658
rect 74454 69606 74466 69658
rect 74518 69606 74540 69658
rect 74188 68570 74540 69606
rect 74188 68518 74210 68570
rect 74262 68518 74274 68570
rect 74326 68518 74338 68570
rect 74390 68518 74402 68570
rect 74454 68518 74466 68570
rect 74518 68518 74540 68570
rect 74188 67482 74540 68518
rect 74188 67430 74210 67482
rect 74262 67430 74274 67482
rect 74326 67430 74338 67482
rect 74390 67430 74402 67482
rect 74454 67430 74466 67482
rect 74518 67430 74540 67482
rect 74188 66394 74540 67430
rect 74188 66342 74210 66394
rect 74262 66342 74274 66394
rect 74326 66342 74338 66394
rect 74390 66342 74402 66394
rect 74454 66342 74466 66394
rect 74518 66342 74540 66394
rect 74188 65306 74540 66342
rect 74188 65254 74210 65306
rect 74262 65254 74274 65306
rect 74326 65254 74338 65306
rect 74390 65254 74402 65306
rect 74454 65254 74466 65306
rect 74518 65254 74540 65306
rect 74188 64588 74540 65254
rect 74188 64532 74216 64588
rect 74272 64532 74296 64588
rect 74352 64532 74376 64588
rect 74432 64532 74456 64588
rect 74512 64532 74540 64588
rect 74188 64508 74540 64532
rect 74188 64452 74216 64508
rect 74272 64452 74296 64508
rect 74352 64452 74376 64508
rect 74432 64452 74456 64508
rect 74512 64452 74540 64508
rect 74188 64428 74540 64452
rect 74188 64372 74216 64428
rect 74272 64372 74296 64428
rect 74352 64372 74376 64428
rect 74432 64372 74456 64428
rect 74512 64372 74540 64428
rect 74188 64348 74540 64372
rect 74188 64292 74216 64348
rect 74272 64292 74296 64348
rect 74352 64292 74376 64348
rect 74432 64292 74456 64348
rect 74512 64292 74540 64348
rect 74188 64218 74540 64292
rect 74188 64166 74210 64218
rect 74262 64166 74274 64218
rect 74326 64166 74338 64218
rect 74390 64166 74402 64218
rect 74454 64166 74466 64218
rect 74518 64166 74540 64218
rect 74188 63130 74540 64166
rect 74188 63078 74210 63130
rect 74262 63078 74274 63130
rect 74326 63078 74338 63130
rect 74390 63078 74402 63130
rect 74454 63078 74466 63130
rect 74518 63078 74540 63130
rect 74188 62042 74540 63078
rect 74188 61990 74210 62042
rect 74262 61990 74274 62042
rect 74326 61990 74338 62042
rect 74390 61990 74402 62042
rect 74454 61990 74466 62042
rect 74518 61990 74540 62042
rect 74188 60954 74540 61990
rect 74188 60902 74210 60954
rect 74262 60902 74274 60954
rect 74326 60902 74338 60954
rect 74390 60902 74402 60954
rect 74454 60902 74466 60954
rect 74518 60902 74540 60954
rect 74188 59866 74540 60902
rect 74188 59814 74210 59866
rect 74262 59814 74274 59866
rect 74326 59814 74338 59866
rect 74390 59814 74402 59866
rect 74454 59814 74466 59866
rect 74518 59814 74540 59866
rect 74188 58778 74540 59814
rect 74188 58726 74210 58778
rect 74262 58726 74274 58778
rect 74326 58726 74338 58778
rect 74390 58726 74402 58778
rect 74454 58726 74466 58778
rect 74518 58726 74540 58778
rect 74188 57690 74540 58726
rect 74188 57638 74210 57690
rect 74262 57638 74274 57690
rect 74326 57638 74338 57690
rect 74390 57638 74402 57690
rect 74454 57638 74466 57690
rect 74518 57638 74540 57690
rect 74188 56602 74540 57638
rect 74188 56550 74210 56602
rect 74262 56550 74274 56602
rect 74326 56550 74338 56602
rect 74390 56550 74402 56602
rect 74454 56550 74466 56602
rect 74518 56550 74540 56602
rect 74188 55514 74540 56550
rect 74188 55462 74210 55514
rect 74262 55462 74274 55514
rect 74326 55462 74338 55514
rect 74390 55462 74402 55514
rect 74454 55462 74466 55514
rect 74518 55462 74540 55514
rect 74188 54588 74540 55462
rect 74188 54532 74216 54588
rect 74272 54532 74296 54588
rect 74352 54532 74376 54588
rect 74432 54532 74456 54588
rect 74512 54532 74540 54588
rect 74188 54508 74540 54532
rect 74188 54452 74216 54508
rect 74272 54452 74296 54508
rect 74352 54452 74376 54508
rect 74432 54452 74456 54508
rect 74512 54452 74540 54508
rect 74188 54428 74540 54452
rect 74188 54426 74216 54428
rect 74272 54426 74296 54428
rect 74352 54426 74376 54428
rect 74432 54426 74456 54428
rect 74512 54426 74540 54428
rect 74188 54374 74210 54426
rect 74272 54374 74274 54426
rect 74454 54374 74456 54426
rect 74518 54374 74540 54426
rect 74188 54372 74216 54374
rect 74272 54372 74296 54374
rect 74352 54372 74376 54374
rect 74432 54372 74456 54374
rect 74512 54372 74540 54374
rect 74188 54348 74540 54372
rect 74188 54292 74216 54348
rect 74272 54292 74296 54348
rect 74352 54292 74376 54348
rect 74432 54292 74456 54348
rect 74512 54292 74540 54348
rect 74188 53338 74540 54292
rect 74188 53286 74210 53338
rect 74262 53286 74274 53338
rect 74326 53286 74338 53338
rect 74390 53286 74402 53338
rect 74454 53286 74466 53338
rect 74518 53286 74540 53338
rect 74188 52250 74540 53286
rect 74188 52198 74210 52250
rect 74262 52198 74274 52250
rect 74326 52198 74338 52250
rect 74390 52198 74402 52250
rect 74454 52198 74466 52250
rect 74518 52198 74540 52250
rect 74188 51162 74540 52198
rect 74188 51110 74210 51162
rect 74262 51110 74274 51162
rect 74326 51110 74338 51162
rect 74390 51110 74402 51162
rect 74454 51110 74466 51162
rect 74518 51110 74540 51162
rect 74188 50074 74540 51110
rect 74188 50022 74210 50074
rect 74262 50022 74274 50074
rect 74326 50022 74338 50074
rect 74390 50022 74402 50074
rect 74454 50022 74466 50074
rect 74518 50022 74540 50074
rect 74188 48986 74540 50022
rect 74188 48934 74210 48986
rect 74262 48934 74274 48986
rect 74326 48934 74338 48986
rect 74390 48934 74402 48986
rect 74454 48934 74466 48986
rect 74518 48934 74540 48986
rect 74188 47898 74540 48934
rect 74188 47846 74210 47898
rect 74262 47846 74274 47898
rect 74326 47846 74338 47898
rect 74390 47846 74402 47898
rect 74454 47846 74466 47898
rect 74518 47846 74540 47898
rect 74188 46810 74540 47846
rect 74188 46758 74210 46810
rect 74262 46758 74274 46810
rect 74326 46758 74338 46810
rect 74390 46758 74402 46810
rect 74454 46758 74466 46810
rect 74518 46758 74540 46810
rect 74188 45722 74540 46758
rect 74188 45670 74210 45722
rect 74262 45670 74274 45722
rect 74326 45670 74338 45722
rect 74390 45670 74402 45722
rect 74454 45670 74466 45722
rect 74518 45670 74540 45722
rect 74188 44634 74540 45670
rect 74188 44582 74210 44634
rect 74262 44588 74274 44634
rect 74326 44588 74338 44634
rect 74390 44588 74402 44634
rect 74454 44588 74466 44634
rect 74272 44582 74274 44588
rect 74454 44582 74456 44588
rect 74518 44582 74540 44634
rect 74188 44532 74216 44582
rect 74272 44532 74296 44582
rect 74352 44532 74376 44582
rect 74432 44532 74456 44582
rect 74512 44532 74540 44582
rect 74188 44508 74540 44532
rect 74188 44452 74216 44508
rect 74272 44452 74296 44508
rect 74352 44452 74376 44508
rect 74432 44452 74456 44508
rect 74512 44452 74540 44508
rect 74188 44428 74540 44452
rect 74188 44372 74216 44428
rect 74272 44372 74296 44428
rect 74352 44372 74376 44428
rect 74432 44372 74456 44428
rect 74512 44372 74540 44428
rect 74188 44348 74540 44372
rect 74188 44292 74216 44348
rect 74272 44292 74296 44348
rect 74352 44292 74376 44348
rect 74432 44292 74456 44348
rect 74512 44292 74540 44348
rect 74188 43546 74540 44292
rect 74188 43494 74210 43546
rect 74262 43494 74274 43546
rect 74326 43494 74338 43546
rect 74390 43494 74402 43546
rect 74454 43494 74466 43546
rect 74518 43494 74540 43546
rect 74188 42458 74540 43494
rect 74188 42406 74210 42458
rect 74262 42406 74274 42458
rect 74326 42406 74338 42458
rect 74390 42406 74402 42458
rect 74454 42406 74466 42458
rect 74518 42406 74540 42458
rect 74188 41370 74540 42406
rect 74188 41318 74210 41370
rect 74262 41318 74274 41370
rect 74326 41318 74338 41370
rect 74390 41318 74402 41370
rect 74454 41318 74466 41370
rect 74518 41318 74540 41370
rect 74188 40282 74540 41318
rect 74188 40230 74210 40282
rect 74262 40230 74274 40282
rect 74326 40230 74338 40282
rect 74390 40230 74402 40282
rect 74454 40230 74466 40282
rect 74518 40230 74540 40282
rect 74188 39194 74540 40230
rect 74188 39142 74210 39194
rect 74262 39142 74274 39194
rect 74326 39142 74338 39194
rect 74390 39142 74402 39194
rect 74454 39142 74466 39194
rect 74518 39142 74540 39194
rect 74188 38106 74540 39142
rect 74188 38054 74210 38106
rect 74262 38054 74274 38106
rect 74326 38054 74338 38106
rect 74390 38054 74402 38106
rect 74454 38054 74466 38106
rect 74518 38054 74540 38106
rect 74188 37018 74540 38054
rect 74188 36966 74210 37018
rect 74262 36966 74274 37018
rect 74326 36966 74338 37018
rect 74390 36966 74402 37018
rect 74454 36966 74466 37018
rect 74518 36966 74540 37018
rect 74188 35930 74540 36966
rect 74188 35878 74210 35930
rect 74262 35878 74274 35930
rect 74326 35878 74338 35930
rect 74390 35878 74402 35930
rect 74454 35878 74466 35930
rect 74518 35878 74540 35930
rect 74188 34842 74540 35878
rect 74188 34790 74210 34842
rect 74262 34790 74274 34842
rect 74326 34790 74338 34842
rect 74390 34790 74402 34842
rect 74454 34790 74466 34842
rect 74518 34790 74540 34842
rect 74188 34588 74540 34790
rect 74188 34532 74216 34588
rect 74272 34532 74296 34588
rect 74352 34532 74376 34588
rect 74432 34532 74456 34588
rect 74512 34532 74540 34588
rect 74188 34508 74540 34532
rect 74188 34452 74216 34508
rect 74272 34452 74296 34508
rect 74352 34452 74376 34508
rect 74432 34452 74456 34508
rect 74512 34452 74540 34508
rect 74188 34428 74540 34452
rect 74188 34372 74216 34428
rect 74272 34372 74296 34428
rect 74352 34372 74376 34428
rect 74432 34372 74456 34428
rect 74512 34372 74540 34428
rect 74188 34348 74540 34372
rect 74188 34292 74216 34348
rect 74272 34292 74296 34348
rect 74352 34292 74376 34348
rect 74432 34292 74456 34348
rect 74512 34292 74540 34348
rect 74188 33754 74540 34292
rect 74188 33702 74210 33754
rect 74262 33702 74274 33754
rect 74326 33702 74338 33754
rect 74390 33702 74402 33754
rect 74454 33702 74466 33754
rect 74518 33702 74540 33754
rect 74188 32666 74540 33702
rect 74188 32614 74210 32666
rect 74262 32614 74274 32666
rect 74326 32614 74338 32666
rect 74390 32614 74402 32666
rect 74454 32614 74466 32666
rect 74518 32614 74540 32666
rect 74188 31578 74540 32614
rect 74188 31526 74210 31578
rect 74262 31526 74274 31578
rect 74326 31526 74338 31578
rect 74390 31526 74402 31578
rect 74454 31526 74466 31578
rect 74518 31526 74540 31578
rect 74188 30490 74540 31526
rect 74188 30438 74210 30490
rect 74262 30438 74274 30490
rect 74326 30438 74338 30490
rect 74390 30438 74402 30490
rect 74454 30438 74466 30490
rect 74518 30438 74540 30490
rect 74188 29402 74540 30438
rect 74188 29350 74210 29402
rect 74262 29350 74274 29402
rect 74326 29350 74338 29402
rect 74390 29350 74402 29402
rect 74454 29350 74466 29402
rect 74518 29350 74540 29402
rect 74188 28314 74540 29350
rect 74188 28262 74210 28314
rect 74262 28262 74274 28314
rect 74326 28262 74338 28314
rect 74390 28262 74402 28314
rect 74454 28262 74466 28314
rect 74518 28262 74540 28314
rect 74188 27226 74540 28262
rect 74188 27174 74210 27226
rect 74262 27174 74274 27226
rect 74326 27174 74338 27226
rect 74390 27174 74402 27226
rect 74454 27174 74466 27226
rect 74518 27174 74540 27226
rect 74188 26138 74540 27174
rect 74188 26086 74210 26138
rect 74262 26086 74274 26138
rect 74326 26086 74338 26138
rect 74390 26086 74402 26138
rect 74454 26086 74466 26138
rect 74518 26086 74540 26138
rect 74188 25050 74540 26086
rect 74188 24998 74210 25050
rect 74262 24998 74274 25050
rect 74326 24998 74338 25050
rect 74390 24998 74402 25050
rect 74454 24998 74466 25050
rect 74518 24998 74540 25050
rect 74188 24588 74540 24998
rect 74188 24532 74216 24588
rect 74272 24532 74296 24588
rect 74352 24532 74376 24588
rect 74432 24532 74456 24588
rect 74512 24532 74540 24588
rect 74188 24508 74540 24532
rect 74188 24452 74216 24508
rect 74272 24452 74296 24508
rect 74352 24452 74376 24508
rect 74432 24452 74456 24508
rect 74512 24452 74540 24508
rect 74188 24428 74540 24452
rect 74188 24372 74216 24428
rect 74272 24372 74296 24428
rect 74352 24372 74376 24428
rect 74432 24372 74456 24428
rect 74512 24372 74540 24428
rect 74188 24348 74540 24372
rect 74188 24292 74216 24348
rect 74272 24292 74296 24348
rect 74352 24292 74376 24348
rect 74432 24292 74456 24348
rect 74512 24292 74540 24348
rect 74188 23962 74540 24292
rect 74188 23910 74210 23962
rect 74262 23910 74274 23962
rect 74326 23910 74338 23962
rect 74390 23910 74402 23962
rect 74454 23910 74466 23962
rect 74518 23910 74540 23962
rect 74188 22874 74540 23910
rect 74188 22822 74210 22874
rect 74262 22822 74274 22874
rect 74326 22822 74338 22874
rect 74390 22822 74402 22874
rect 74454 22822 74466 22874
rect 74518 22822 74540 22874
rect 74188 21786 74540 22822
rect 74188 21734 74210 21786
rect 74262 21734 74274 21786
rect 74326 21734 74338 21786
rect 74390 21734 74402 21786
rect 74454 21734 74466 21786
rect 74518 21734 74540 21786
rect 74188 20698 74540 21734
rect 74188 20646 74210 20698
rect 74262 20646 74274 20698
rect 74326 20646 74338 20698
rect 74390 20646 74402 20698
rect 74454 20646 74466 20698
rect 74518 20646 74540 20698
rect 74188 19610 74540 20646
rect 74188 19558 74210 19610
rect 74262 19558 74274 19610
rect 74326 19558 74338 19610
rect 74390 19558 74402 19610
rect 74454 19558 74466 19610
rect 74518 19558 74540 19610
rect 74188 18522 74540 19558
rect 74188 18470 74210 18522
rect 74262 18470 74274 18522
rect 74326 18470 74338 18522
rect 74390 18470 74402 18522
rect 74454 18470 74466 18522
rect 74518 18470 74540 18522
rect 74188 17434 74540 18470
rect 74188 17382 74210 17434
rect 74262 17382 74274 17434
rect 74326 17382 74338 17434
rect 74390 17382 74402 17434
rect 74454 17382 74466 17434
rect 74518 17382 74540 17434
rect 74188 16346 74540 17382
rect 74188 16294 74210 16346
rect 74262 16294 74274 16346
rect 74326 16294 74338 16346
rect 74390 16294 74402 16346
rect 74454 16294 74466 16346
rect 74518 16294 74540 16346
rect 74188 15258 74540 16294
rect 74188 15206 74210 15258
rect 74262 15206 74274 15258
rect 74326 15206 74338 15258
rect 74390 15206 74402 15258
rect 74454 15206 74466 15258
rect 74518 15206 74540 15258
rect 74188 14588 74540 15206
rect 74188 14532 74216 14588
rect 74272 14532 74296 14588
rect 74352 14532 74376 14588
rect 74432 14532 74456 14588
rect 74512 14532 74540 14588
rect 74188 14508 74540 14532
rect 74188 14452 74216 14508
rect 74272 14452 74296 14508
rect 74352 14452 74376 14508
rect 74432 14452 74456 14508
rect 74512 14452 74540 14508
rect 74188 14428 74540 14452
rect 74188 14372 74216 14428
rect 74272 14372 74296 14428
rect 74352 14372 74376 14428
rect 74432 14372 74456 14428
rect 74512 14372 74540 14428
rect 74188 14348 74540 14372
rect 74188 14292 74216 14348
rect 74272 14292 74296 14348
rect 74352 14292 74376 14348
rect 74432 14292 74456 14348
rect 74512 14292 74540 14348
rect 74188 14170 74540 14292
rect 74188 14118 74210 14170
rect 74262 14118 74274 14170
rect 74326 14118 74338 14170
rect 74390 14118 74402 14170
rect 74454 14118 74466 14170
rect 74518 14118 74540 14170
rect 74188 13082 74540 14118
rect 74188 13030 74210 13082
rect 74262 13030 74274 13082
rect 74326 13030 74338 13082
rect 74390 13030 74402 13082
rect 74454 13030 74466 13082
rect 74518 13030 74540 13082
rect 74188 11994 74540 13030
rect 74188 11942 74210 11994
rect 74262 11942 74274 11994
rect 74326 11942 74338 11994
rect 74390 11942 74402 11994
rect 74454 11942 74466 11994
rect 74518 11942 74540 11994
rect 74188 10906 74540 11942
rect 74188 10854 74210 10906
rect 74262 10854 74274 10906
rect 74326 10854 74338 10906
rect 74390 10854 74402 10906
rect 74454 10854 74466 10906
rect 74518 10854 74540 10906
rect 74188 9818 74540 10854
rect 74188 9766 74210 9818
rect 74262 9766 74274 9818
rect 74326 9766 74338 9818
rect 74390 9766 74402 9818
rect 74454 9766 74466 9818
rect 74518 9766 74540 9818
rect 74188 8730 74540 9766
rect 74188 8678 74210 8730
rect 74262 8678 74274 8730
rect 74326 8678 74338 8730
rect 74390 8678 74402 8730
rect 74454 8678 74466 8730
rect 74518 8678 74540 8730
rect 74188 7642 74540 8678
rect 74188 7590 74210 7642
rect 74262 7590 74274 7642
rect 74326 7590 74338 7642
rect 74390 7590 74402 7642
rect 74454 7590 74466 7642
rect 74518 7590 74540 7642
rect 74188 6554 74540 7590
rect 74188 6502 74210 6554
rect 74262 6502 74274 6554
rect 74326 6502 74338 6554
rect 74390 6502 74402 6554
rect 74454 6502 74466 6554
rect 74518 6502 74540 6554
rect 74188 5466 74540 6502
rect 74188 5414 74210 5466
rect 74262 5414 74274 5466
rect 74326 5414 74338 5466
rect 74390 5414 74402 5466
rect 74454 5414 74466 5466
rect 74518 5414 74540 5466
rect 74188 4588 74540 5414
rect 74188 4532 74216 4588
rect 74272 4532 74296 4588
rect 74352 4532 74376 4588
rect 74432 4532 74456 4588
rect 74512 4532 74540 4588
rect 74188 4508 74540 4532
rect 74188 4452 74216 4508
rect 74272 4452 74296 4508
rect 74352 4452 74376 4508
rect 74432 4452 74456 4508
rect 74512 4452 74540 4508
rect 74188 4428 74540 4452
rect 74188 4378 74216 4428
rect 74272 4378 74296 4428
rect 74352 4378 74376 4428
rect 74432 4378 74456 4428
rect 74512 4378 74540 4428
rect 74188 4326 74210 4378
rect 74272 4372 74274 4378
rect 74454 4372 74456 4378
rect 74262 4348 74274 4372
rect 74326 4348 74338 4372
rect 74390 4348 74402 4372
rect 74454 4348 74466 4372
rect 74272 4326 74274 4348
rect 74454 4326 74456 4348
rect 74518 4326 74540 4378
rect 74188 4292 74216 4326
rect 74272 4292 74296 4326
rect 74352 4292 74376 4326
rect 74432 4292 74456 4326
rect 74512 4292 74540 4326
rect 74188 3290 74540 4292
rect 74188 3238 74210 3290
rect 74262 3238 74274 3290
rect 74326 3238 74338 3290
rect 74390 3238 74402 3290
rect 74454 3238 74466 3290
rect 74518 3238 74540 3290
rect 72608 2440 72660 2446
rect 72608 2382 72660 2388
rect 71836 2180 71864 2236
rect 71920 2180 71944 2236
rect 72000 2180 72024 2236
rect 72080 2180 72104 2236
rect 72160 2180 72188 2236
rect 71836 2156 72188 2180
rect 71836 2100 71864 2156
rect 71920 2100 71944 2156
rect 72000 2100 72024 2156
rect 72080 2100 72104 2156
rect 72160 2100 72188 2156
rect 71836 2076 72188 2100
rect 71836 2020 71864 2076
rect 71920 2020 71944 2076
rect 72000 2020 72024 2076
rect 72080 2020 72104 2076
rect 72160 2020 72188 2076
rect 71836 1996 72188 2020
rect 70860 1964 70912 1970
rect 70860 1906 70912 1912
rect 71412 1964 71464 1970
rect 71412 1906 71464 1912
rect 71836 1940 71864 1996
rect 71920 1940 71944 1996
rect 72000 1940 72024 1996
rect 72080 1940 72104 1996
rect 72160 1940 72188 1996
rect 71320 1896 71372 1902
rect 71320 1838 71372 1844
rect 70584 1352 70636 1358
rect 70584 1294 70636 1300
rect 70860 1352 70912 1358
rect 70860 1294 70912 1300
rect 70872 800 70900 1294
rect 71332 800 71360 1838
rect 71836 1658 72188 1940
rect 71836 1606 71858 1658
rect 71910 1606 71922 1658
rect 71974 1606 71986 1658
rect 72038 1606 72050 1658
rect 72102 1606 72114 1658
rect 72166 1606 72188 1658
rect 71836 1040 72188 1606
rect 72620 1290 72648 2382
rect 74188 2202 74540 3238
rect 74188 2150 74210 2202
rect 74262 2150 74274 2202
rect 74326 2150 74338 2202
rect 74390 2150 74402 2202
rect 74454 2150 74466 2202
rect 74518 2150 74540 2202
rect 72608 1284 72660 1290
rect 72608 1226 72660 1232
rect 74188 1114 74540 2150
rect 74188 1062 74210 1114
rect 74262 1062 74274 1114
rect 74326 1062 74338 1114
rect 74390 1062 74402 1114
rect 74454 1062 74466 1114
rect 74518 1062 74540 1114
rect 74188 1040 74540 1062
rect 65708 128 65760 134
rect 65708 70 65760 76
rect 65798 0 65854 800
rect 66258 0 66314 800
rect 66718 0 66774 800
rect 67178 0 67234 800
rect 67638 0 67694 800
rect 68098 0 68154 800
rect 68558 0 68614 800
rect 69018 0 69074 800
rect 69478 0 69534 800
rect 69938 0 69994 800
rect 70398 0 70454 800
rect 70858 0 70914 800
rect 71318 0 71374 800
<< via2 >>
rect 2136 84532 2192 84588
rect 2136 84452 2192 84508
rect 2136 84372 2192 84428
rect 2136 84292 2192 84348
rect 5632 84532 5688 84588
rect 5632 84452 5688 84508
rect 5632 84372 5688 84428
rect 5632 84292 5688 84348
rect 8522 84532 8578 84588
rect 8522 84452 8578 84508
rect 8522 84372 8578 84428
rect 8522 84292 8578 84348
rect 11412 84532 11468 84588
rect 11412 84452 11468 84508
rect 11412 84372 11468 84428
rect 11412 84292 11468 84348
rect 14302 84532 14358 84588
rect 14302 84452 14358 84508
rect 14302 84372 14358 84428
rect 14302 84292 14358 84348
rect 17192 84532 17248 84588
rect 17192 84452 17248 84508
rect 17192 84372 17248 84428
rect 17192 84292 17248 84348
rect 20082 84532 20138 84588
rect 20082 84452 20138 84508
rect 20082 84372 20138 84428
rect 20082 84292 20138 84348
rect 22972 84532 23028 84588
rect 22972 84452 23028 84508
rect 22972 84372 23028 84428
rect 22972 84292 23028 84348
rect 25862 84532 25918 84588
rect 25862 84452 25918 84508
rect 25862 84372 25918 84428
rect 25862 84292 25918 84348
rect 28752 84532 28808 84588
rect 28752 84452 28808 84508
rect 28752 84372 28808 84428
rect 28752 84292 28808 84348
rect 31642 84532 31698 84588
rect 31642 84452 31698 84508
rect 31642 84372 31698 84428
rect 31642 84292 31698 84348
rect 34532 84532 34588 84588
rect 34532 84452 34588 84508
rect 34532 84372 34588 84428
rect 34532 84292 34588 84348
rect 37422 84532 37478 84588
rect 37422 84452 37478 84508
rect 37422 84372 37478 84428
rect 37422 84292 37478 84348
rect 40312 84532 40368 84588
rect 40312 84452 40368 84508
rect 40312 84372 40368 84428
rect 40312 84292 40368 84348
rect 43202 84532 43258 84588
rect 43202 84452 43258 84508
rect 43202 84372 43258 84428
rect 43202 84292 43258 84348
rect 46092 84532 46148 84588
rect 46092 84452 46148 84508
rect 46092 84372 46148 84428
rect 46092 84292 46148 84348
rect 49100 84532 49156 84588
rect 49100 84452 49156 84508
rect 49100 84372 49156 84428
rect 49100 84292 49156 84348
rect 52329 84532 52385 84588
rect 52329 84452 52385 84508
rect 52329 84372 52385 84428
rect 52329 84292 52385 84348
rect 53730 84532 53786 84588
rect 53730 84452 53786 84508
rect 53730 84372 53786 84428
rect 53730 84292 53786 84348
rect 53898 84532 53954 84588
rect 53898 84452 53954 84508
rect 53898 84372 53954 84428
rect 53898 84292 53954 84348
rect 54642 84532 54698 84588
rect 54642 84452 54698 84508
rect 54642 84372 54698 84428
rect 54642 84292 54698 84348
rect 55032 84532 55088 84588
rect 55032 84452 55088 84508
rect 55032 84372 55088 84428
rect 55032 84292 55088 84348
rect 55748 84532 55804 84588
rect 55748 84452 55804 84508
rect 55748 84372 55804 84428
rect 55748 84292 55804 84348
rect 56326 84532 56382 84588
rect 56326 84452 56382 84508
rect 56326 84372 56382 84428
rect 56326 84292 56382 84348
rect 56771 84532 56827 84588
rect 56771 84452 56827 84508
rect 56771 84372 56827 84428
rect 56771 84292 56827 84348
rect 57075 84532 57131 84588
rect 57075 84452 57131 84508
rect 57075 84372 57131 84428
rect 57075 84292 57131 84348
rect 57917 84532 57973 84588
rect 57917 84452 57973 84508
rect 57917 84372 57973 84428
rect 57917 84292 57973 84348
rect 58557 84532 58613 84588
rect 58557 84452 58613 84508
rect 58557 84372 58613 84428
rect 58557 84292 58613 84348
rect 59140 84532 59196 84588
rect 59140 84452 59196 84508
rect 59140 84372 59196 84428
rect 59140 84292 59196 84348
rect 60418 84532 60474 84588
rect 60418 84452 60474 84508
rect 60418 84372 60474 84428
rect 60418 84292 60474 84348
rect 60576 84532 60632 84588
rect 60576 84452 60632 84508
rect 60576 84372 60632 84428
rect 60576 84292 60632 84348
rect 62620 84532 62676 84588
rect 62700 84532 62756 84588
rect 62620 84452 62676 84508
rect 62700 84452 62756 84508
rect 62620 84372 62676 84428
rect 62700 84372 62756 84428
rect 62620 84292 62676 84348
rect 62700 84292 62756 84348
rect 2276 82180 2332 82236
rect 2356 82180 2412 82236
rect 2276 82100 2332 82156
rect 2356 82100 2412 82156
rect 2276 82020 2332 82076
rect 2356 82020 2412 82076
rect 2276 81940 2332 81996
rect 2356 81940 2412 81996
rect 5485 82180 5541 82236
rect 5485 82100 5541 82156
rect 5485 82020 5541 82076
rect 5485 81940 5541 81996
rect 8375 82180 8431 82236
rect 8375 82100 8431 82156
rect 8375 82020 8431 82076
rect 8375 81940 8431 81996
rect 11265 82180 11321 82236
rect 11265 82100 11321 82156
rect 11265 82020 11321 82076
rect 11265 81940 11321 81996
rect 14155 82180 14211 82236
rect 14155 82100 14211 82156
rect 14155 82020 14211 82076
rect 14155 81940 14211 81996
rect 17045 82180 17101 82236
rect 17045 82100 17101 82156
rect 17045 82020 17101 82076
rect 17045 81940 17101 81996
rect 19935 82180 19991 82236
rect 19935 82100 19991 82156
rect 19935 82020 19991 82076
rect 19935 81940 19991 81996
rect 22825 82180 22881 82236
rect 22825 82100 22881 82156
rect 22825 82020 22881 82076
rect 22825 81940 22881 81996
rect 25715 82180 25771 82236
rect 25715 82100 25771 82156
rect 25715 82020 25771 82076
rect 25715 81940 25771 81996
rect 28605 82180 28661 82236
rect 28605 82100 28661 82156
rect 28605 82020 28661 82076
rect 28605 81940 28661 81996
rect 31495 82180 31551 82236
rect 31495 82100 31551 82156
rect 31495 82020 31551 82076
rect 31495 81940 31551 81996
rect 34385 82180 34441 82236
rect 34385 82100 34441 82156
rect 34385 82020 34441 82076
rect 34385 81940 34441 81996
rect 37275 82180 37331 82236
rect 37275 82100 37331 82156
rect 37275 82020 37331 82076
rect 37275 81940 37331 81996
rect 40165 82180 40221 82236
rect 40165 82100 40221 82156
rect 40165 82020 40221 82076
rect 40165 81940 40221 81996
rect 43055 82180 43111 82236
rect 43055 82100 43111 82156
rect 43055 82020 43111 82076
rect 43055 81940 43111 81996
rect 45945 82180 46001 82236
rect 45945 82100 46001 82156
rect 45945 82020 46001 82076
rect 45945 81940 46001 81996
rect 48892 82180 48948 82236
rect 48892 82100 48948 82156
rect 48892 82020 48948 82076
rect 48892 81940 48948 81996
rect 49754 82180 49810 82236
rect 49834 82180 49890 82236
rect 49754 82100 49810 82156
rect 49834 82100 49890 82156
rect 49754 82020 49810 82076
rect 49834 82020 49890 82076
rect 49754 81940 49810 81996
rect 49834 81940 49890 81996
rect 53048 82180 53104 82236
rect 53048 82100 53104 82156
rect 53048 82020 53104 82076
rect 53048 81940 53104 81996
rect 53206 82180 53262 82236
rect 53206 82100 53262 82156
rect 53206 82020 53262 82076
rect 53206 81940 53262 81996
rect 53562 82180 53618 82236
rect 53562 82100 53618 82156
rect 53562 82020 53618 82076
rect 53562 81940 53618 81996
rect 54880 82180 54936 82236
rect 54880 82100 54936 82156
rect 54880 82020 54936 82076
rect 54880 81940 54936 81996
rect 55473 82180 55529 82236
rect 55473 82100 55529 82156
rect 55473 82020 55529 82076
rect 55473 81940 55529 81996
rect 56619 82180 56675 82236
rect 56619 82100 56675 82156
rect 56619 82020 56675 82076
rect 56619 81940 56675 81996
rect 58055 82180 58111 82236
rect 58135 82180 58191 82236
rect 58055 82100 58111 82156
rect 58135 82100 58191 82156
rect 58055 82020 58111 82076
rect 58135 82020 58191 82076
rect 58055 81940 58111 81996
rect 58135 81940 58191 81996
rect 59298 82180 59354 82236
rect 59298 82100 59354 82156
rect 59298 82020 59354 82076
rect 59298 81940 59354 81996
rect 59456 82180 59512 82236
rect 59456 82100 59512 82156
rect 59456 82020 59512 82076
rect 59456 81940 59512 81996
rect 59764 82180 59820 82236
rect 59764 82100 59820 82156
rect 59764 82020 59820 82076
rect 59764 81940 59820 81996
rect 59910 82180 59966 82236
rect 59910 82100 59966 82156
rect 59910 82020 59966 82076
rect 59910 81940 59966 81996
rect 60046 82180 60102 82236
rect 60126 82180 60182 82236
rect 60046 82100 60102 82156
rect 60126 82100 60182 82156
rect 60046 82020 60102 82076
rect 60126 82020 60182 82076
rect 60046 81940 60102 81996
rect 60126 81940 60182 81996
rect 62418 82180 62474 82236
rect 62498 82180 62554 82236
rect 62418 82100 62474 82156
rect 62498 82100 62554 82156
rect 62418 82020 62474 82076
rect 62498 82020 62554 82076
rect 62418 81940 62474 81996
rect 62498 81940 62554 81996
rect 2136 74532 2192 74588
rect 2136 74452 2192 74508
rect 2136 74372 2192 74428
rect 2136 74292 2192 74348
rect 5632 74532 5688 74588
rect 5632 74452 5688 74508
rect 5632 74372 5688 74428
rect 5632 74292 5688 74348
rect 8522 74532 8578 74588
rect 8522 74452 8578 74508
rect 8522 74372 8578 74428
rect 8522 74292 8578 74348
rect 11412 74532 11468 74588
rect 11412 74452 11468 74508
rect 11412 74372 11468 74428
rect 11412 74292 11468 74348
rect 14302 74532 14358 74588
rect 14302 74452 14358 74508
rect 14302 74372 14358 74428
rect 14302 74292 14358 74348
rect 17192 74532 17248 74588
rect 17192 74452 17248 74508
rect 17192 74372 17248 74428
rect 17192 74292 17248 74348
rect 20082 74532 20138 74588
rect 20082 74452 20138 74508
rect 20082 74372 20138 74428
rect 20082 74292 20138 74348
rect 22972 74532 23028 74588
rect 22972 74452 23028 74508
rect 22972 74372 23028 74428
rect 22972 74292 23028 74348
rect 25862 74532 25918 74588
rect 25862 74452 25918 74508
rect 25862 74372 25918 74428
rect 25862 74292 25918 74348
rect 28752 74532 28808 74588
rect 28752 74452 28808 74508
rect 28752 74372 28808 74428
rect 28752 74292 28808 74348
rect 31642 74532 31698 74588
rect 31642 74452 31698 74508
rect 31642 74372 31698 74428
rect 31642 74292 31698 74348
rect 34532 74532 34588 74588
rect 34532 74452 34588 74508
rect 34532 74372 34588 74428
rect 34532 74292 34588 74348
rect 37422 74532 37478 74588
rect 37422 74452 37478 74508
rect 37422 74372 37478 74428
rect 37422 74292 37478 74348
rect 40312 74532 40368 74588
rect 40312 74452 40368 74508
rect 40312 74372 40368 74428
rect 40312 74292 40368 74348
rect 43202 74532 43258 74588
rect 43202 74452 43258 74508
rect 43202 74372 43258 74428
rect 43202 74292 43258 74348
rect 46092 74532 46148 74588
rect 46092 74452 46148 74508
rect 46092 74372 46148 74428
rect 46092 74292 46148 74348
rect 49100 74532 49156 74588
rect 49100 74452 49156 74508
rect 49100 74372 49156 74428
rect 49100 74292 49156 74348
rect 52329 74532 52385 74588
rect 52329 74452 52385 74508
rect 52329 74372 52385 74428
rect 52329 74292 52385 74348
rect 53730 74532 53786 74588
rect 53730 74452 53786 74508
rect 53730 74372 53786 74428
rect 53730 74292 53786 74348
rect 53898 74532 53954 74588
rect 53898 74452 53954 74508
rect 53898 74372 53954 74428
rect 53898 74292 53954 74348
rect 54642 74532 54698 74588
rect 54642 74452 54698 74508
rect 54642 74372 54698 74428
rect 54642 74292 54698 74348
rect 55032 74532 55088 74588
rect 55032 74452 55088 74508
rect 55032 74372 55088 74428
rect 55032 74292 55088 74348
rect 55748 74532 55804 74588
rect 55748 74452 55804 74508
rect 55748 74372 55804 74428
rect 55748 74292 55804 74348
rect 56326 74532 56382 74588
rect 56326 74452 56382 74508
rect 56326 74372 56382 74428
rect 56326 74292 56382 74348
rect 56771 74532 56827 74588
rect 56771 74452 56827 74508
rect 56771 74372 56827 74428
rect 56771 74292 56827 74348
rect 57075 74532 57131 74588
rect 57075 74452 57131 74508
rect 57075 74372 57131 74428
rect 57075 74292 57131 74348
rect 57917 74532 57973 74588
rect 57917 74452 57973 74508
rect 57917 74372 57973 74428
rect 57917 74292 57973 74348
rect 58557 74532 58613 74588
rect 58557 74452 58613 74508
rect 58557 74372 58613 74428
rect 58557 74292 58613 74348
rect 59140 74532 59196 74588
rect 59140 74452 59196 74508
rect 59140 74372 59196 74428
rect 59140 74292 59196 74348
rect 60418 74532 60474 74588
rect 60418 74452 60474 74508
rect 60418 74372 60474 74428
rect 60418 74292 60474 74348
rect 60576 74532 60632 74588
rect 60576 74452 60632 74508
rect 60576 74372 60632 74428
rect 60576 74292 60632 74348
rect 62620 74532 62676 74588
rect 62700 74532 62756 74588
rect 62620 74452 62676 74508
rect 62700 74452 62756 74508
rect 62620 74372 62676 74428
rect 62700 74372 62756 74428
rect 62620 74292 62676 74348
rect 62700 74292 62756 74348
rect 2276 72180 2332 72236
rect 2356 72180 2412 72236
rect 2276 72100 2332 72156
rect 2356 72100 2412 72156
rect 2276 72020 2332 72076
rect 2356 72020 2412 72076
rect 2276 71940 2332 71996
rect 2356 71940 2412 71996
rect 5485 72180 5541 72236
rect 5485 72100 5541 72156
rect 5485 72020 5541 72076
rect 5485 71940 5541 71996
rect 8375 72180 8431 72236
rect 8375 72100 8431 72156
rect 8375 72020 8431 72076
rect 8375 71940 8431 71996
rect 11265 72180 11321 72236
rect 11265 72100 11321 72156
rect 11265 72020 11321 72076
rect 11265 71940 11321 71996
rect 14155 72180 14211 72236
rect 14155 72100 14211 72156
rect 14155 72020 14211 72076
rect 14155 71940 14211 71996
rect 17045 72180 17101 72236
rect 17045 72100 17101 72156
rect 17045 72020 17101 72076
rect 17045 71940 17101 71996
rect 19935 72180 19991 72236
rect 19935 72100 19991 72156
rect 19935 72020 19991 72076
rect 19935 71940 19991 71996
rect 22825 72180 22881 72236
rect 22825 72100 22881 72156
rect 22825 72020 22881 72076
rect 22825 71940 22881 71996
rect 25715 72180 25771 72236
rect 25715 72100 25771 72156
rect 25715 72020 25771 72076
rect 25715 71940 25771 71996
rect 28605 72180 28661 72236
rect 28605 72100 28661 72156
rect 28605 72020 28661 72076
rect 28605 71940 28661 71996
rect 31495 72180 31551 72236
rect 31495 72100 31551 72156
rect 31495 72020 31551 72076
rect 31495 71940 31551 71996
rect 34385 72180 34441 72236
rect 34385 72100 34441 72156
rect 34385 72020 34441 72076
rect 34385 71940 34441 71996
rect 37275 72180 37331 72236
rect 37275 72100 37331 72156
rect 37275 72020 37331 72076
rect 37275 71940 37331 71996
rect 40165 72180 40221 72236
rect 40165 72100 40221 72156
rect 40165 72020 40221 72076
rect 40165 71940 40221 71996
rect 43055 72180 43111 72236
rect 43055 72100 43111 72156
rect 43055 72020 43111 72076
rect 43055 71940 43111 71996
rect 45945 72180 46001 72236
rect 45945 72100 46001 72156
rect 45945 72020 46001 72076
rect 45945 71940 46001 71996
rect 48892 72180 48948 72236
rect 48892 72100 48948 72156
rect 48892 72020 48948 72076
rect 48892 71940 48948 71996
rect 49754 72180 49810 72236
rect 49834 72180 49890 72236
rect 49754 72100 49810 72156
rect 49834 72100 49890 72156
rect 49754 72020 49810 72076
rect 49834 72020 49890 72076
rect 49754 71940 49810 71996
rect 49834 71940 49890 71996
rect 53048 72180 53104 72236
rect 53048 72100 53104 72156
rect 53048 72020 53104 72076
rect 53048 71940 53104 71996
rect 53206 72180 53262 72236
rect 53206 72100 53262 72156
rect 53206 72020 53262 72076
rect 53206 71940 53262 71996
rect 53562 72180 53618 72236
rect 53562 72100 53618 72156
rect 53562 72020 53618 72076
rect 53562 71940 53618 71996
rect 54880 72180 54936 72236
rect 54880 72100 54936 72156
rect 54880 72020 54936 72076
rect 54880 71940 54936 71996
rect 55473 72180 55529 72236
rect 55473 72100 55529 72156
rect 55473 72020 55529 72076
rect 55473 71940 55529 71996
rect 56619 72180 56675 72236
rect 56619 72100 56675 72156
rect 56619 72020 56675 72076
rect 56619 71940 56675 71996
rect 58055 72180 58111 72236
rect 58135 72180 58191 72236
rect 58055 72100 58111 72156
rect 58135 72100 58191 72156
rect 58055 72020 58111 72076
rect 58135 72020 58191 72076
rect 58055 71940 58111 71996
rect 58135 71940 58191 71996
rect 59298 72180 59354 72236
rect 59298 72100 59354 72156
rect 59298 72020 59354 72076
rect 59298 71940 59354 71996
rect 59456 72180 59512 72236
rect 59456 72100 59512 72156
rect 59456 72020 59512 72076
rect 59456 71940 59512 71996
rect 59764 72180 59820 72236
rect 59764 72100 59820 72156
rect 59764 72020 59820 72076
rect 59764 71940 59820 71996
rect 59910 72180 59966 72236
rect 59910 72100 59966 72156
rect 59910 72020 59966 72076
rect 59910 71940 59966 71996
rect 60046 72180 60102 72236
rect 60126 72180 60182 72236
rect 60046 72100 60102 72156
rect 60126 72100 60182 72156
rect 60046 72020 60102 72076
rect 60126 72020 60182 72076
rect 60046 71940 60102 71996
rect 60126 71940 60182 71996
rect 62418 72180 62474 72236
rect 62498 72180 62554 72236
rect 62418 72100 62474 72156
rect 62498 72100 62554 72156
rect 62418 72020 62474 72076
rect 62498 72020 62554 72076
rect 62418 71940 62474 71996
rect 62498 71940 62554 71996
rect 63498 65220 63500 65240
rect 63500 65220 63552 65240
rect 63552 65220 63554 65240
rect 63498 65184 63554 65220
rect 2136 64532 2192 64588
rect 2136 64452 2192 64508
rect 2136 64372 2192 64428
rect 2136 64292 2192 64348
rect 5632 64532 5688 64588
rect 5632 64452 5688 64508
rect 5632 64372 5688 64428
rect 5632 64292 5688 64348
rect 8522 64532 8578 64588
rect 8522 64452 8578 64508
rect 8522 64372 8578 64428
rect 8522 64292 8578 64348
rect 11412 64532 11468 64588
rect 11412 64452 11468 64508
rect 11412 64372 11468 64428
rect 11412 64292 11468 64348
rect 14302 64532 14358 64588
rect 14302 64452 14358 64508
rect 14302 64372 14358 64428
rect 14302 64292 14358 64348
rect 17192 64532 17248 64588
rect 17192 64452 17248 64508
rect 17192 64372 17248 64428
rect 17192 64292 17248 64348
rect 20082 64532 20138 64588
rect 20082 64452 20138 64508
rect 20082 64372 20138 64428
rect 20082 64292 20138 64348
rect 22972 64532 23028 64588
rect 22972 64452 23028 64508
rect 22972 64372 23028 64428
rect 22972 64292 23028 64348
rect 25862 64532 25918 64588
rect 25862 64452 25918 64508
rect 25862 64372 25918 64428
rect 25862 64292 25918 64348
rect 28752 64532 28808 64588
rect 28752 64452 28808 64508
rect 28752 64372 28808 64428
rect 28752 64292 28808 64348
rect 31642 64532 31698 64588
rect 31642 64452 31698 64508
rect 31642 64372 31698 64428
rect 31642 64292 31698 64348
rect 34532 64532 34588 64588
rect 34532 64452 34588 64508
rect 34532 64372 34588 64428
rect 34532 64292 34588 64348
rect 37422 64532 37478 64588
rect 37422 64452 37478 64508
rect 37422 64372 37478 64428
rect 37422 64292 37478 64348
rect 40312 64532 40368 64588
rect 40312 64452 40368 64508
rect 40312 64372 40368 64428
rect 40312 64292 40368 64348
rect 43202 64532 43258 64588
rect 43202 64452 43258 64508
rect 43202 64372 43258 64428
rect 43202 64292 43258 64348
rect 46092 64532 46148 64588
rect 46092 64452 46148 64508
rect 46092 64372 46148 64428
rect 46092 64292 46148 64348
rect 49100 64532 49156 64588
rect 49100 64452 49156 64508
rect 49100 64372 49156 64428
rect 49100 64292 49156 64348
rect 52329 64532 52385 64588
rect 52329 64452 52385 64508
rect 52329 64372 52385 64428
rect 52329 64292 52385 64348
rect 53730 64532 53786 64588
rect 53730 64452 53786 64508
rect 53730 64372 53786 64428
rect 53730 64292 53786 64348
rect 53898 64532 53954 64588
rect 53898 64452 53954 64508
rect 53898 64372 53954 64428
rect 53898 64292 53954 64348
rect 54642 64532 54698 64588
rect 54642 64452 54698 64508
rect 54642 64372 54698 64428
rect 54642 64292 54698 64348
rect 55032 64532 55088 64588
rect 55032 64452 55088 64508
rect 55032 64372 55088 64428
rect 55032 64292 55088 64348
rect 55748 64532 55804 64588
rect 55748 64452 55804 64508
rect 55748 64372 55804 64428
rect 55748 64292 55804 64348
rect 56326 64532 56382 64588
rect 56326 64452 56382 64508
rect 56326 64372 56382 64428
rect 56326 64292 56382 64348
rect 56771 64532 56827 64588
rect 56771 64452 56827 64508
rect 56771 64372 56827 64428
rect 56771 64292 56827 64348
rect 57075 64532 57131 64588
rect 57075 64452 57131 64508
rect 57075 64372 57131 64428
rect 57075 64292 57131 64348
rect 57917 64532 57973 64588
rect 57917 64452 57973 64508
rect 57917 64372 57973 64428
rect 57917 64292 57973 64348
rect 58557 64532 58613 64588
rect 58557 64452 58613 64508
rect 58557 64372 58613 64428
rect 58557 64292 58613 64348
rect 59140 64532 59196 64588
rect 59140 64452 59196 64508
rect 59140 64372 59196 64428
rect 59140 64292 59196 64348
rect 60418 64532 60474 64588
rect 60418 64452 60474 64508
rect 60418 64372 60474 64428
rect 60418 64292 60474 64348
rect 60576 64532 60632 64588
rect 60576 64452 60632 64508
rect 60576 64372 60632 64428
rect 60576 64292 60632 64348
rect 62620 64532 62676 64588
rect 62700 64532 62756 64588
rect 62620 64452 62676 64508
rect 62700 64452 62756 64508
rect 62620 64372 62676 64428
rect 62700 64372 62756 64428
rect 62620 64292 62676 64348
rect 62700 64292 62756 64348
rect 63498 63180 63500 63200
rect 63500 63180 63552 63200
rect 63552 63180 63554 63200
rect 63498 63144 63554 63180
rect 2276 62180 2332 62236
rect 2356 62180 2412 62236
rect 2276 62100 2332 62156
rect 2356 62100 2412 62156
rect 2276 62020 2332 62076
rect 2356 62020 2412 62076
rect 2276 61940 2332 61996
rect 2356 61940 2412 61996
rect 5485 62180 5541 62236
rect 5485 62100 5541 62156
rect 5485 62020 5541 62076
rect 5485 61940 5541 61996
rect 8375 62180 8431 62236
rect 8375 62100 8431 62156
rect 8375 62020 8431 62076
rect 8375 61940 8431 61996
rect 11265 62180 11321 62236
rect 11265 62100 11321 62156
rect 11265 62020 11321 62076
rect 11265 61940 11321 61996
rect 14155 62180 14211 62236
rect 14155 62100 14211 62156
rect 14155 62020 14211 62076
rect 14155 61940 14211 61996
rect 17045 62180 17101 62236
rect 17045 62100 17101 62156
rect 17045 62020 17101 62076
rect 17045 61940 17101 61996
rect 19935 62180 19991 62236
rect 19935 62100 19991 62156
rect 19935 62020 19991 62076
rect 19935 61940 19991 61996
rect 22825 62180 22881 62236
rect 22825 62100 22881 62156
rect 22825 62020 22881 62076
rect 22825 61940 22881 61996
rect 25715 62180 25771 62236
rect 25715 62100 25771 62156
rect 25715 62020 25771 62076
rect 25715 61940 25771 61996
rect 28605 62180 28661 62236
rect 28605 62100 28661 62156
rect 28605 62020 28661 62076
rect 28605 61940 28661 61996
rect 31495 62180 31551 62236
rect 31495 62100 31551 62156
rect 31495 62020 31551 62076
rect 31495 61940 31551 61996
rect 34385 62180 34441 62236
rect 34385 62100 34441 62156
rect 34385 62020 34441 62076
rect 34385 61940 34441 61996
rect 37275 62180 37331 62236
rect 37275 62100 37331 62156
rect 37275 62020 37331 62076
rect 37275 61940 37331 61996
rect 40165 62180 40221 62236
rect 40165 62100 40221 62156
rect 40165 62020 40221 62076
rect 40165 61940 40221 61996
rect 43055 62180 43111 62236
rect 43055 62100 43111 62156
rect 43055 62020 43111 62076
rect 43055 61940 43111 61996
rect 45945 62180 46001 62236
rect 45945 62100 46001 62156
rect 45945 62020 46001 62076
rect 45945 61940 46001 61996
rect 48892 62180 48948 62236
rect 48892 62100 48948 62156
rect 48892 62020 48948 62076
rect 48892 61940 48948 61996
rect 49754 62180 49810 62236
rect 49834 62180 49890 62236
rect 49754 62100 49810 62156
rect 49834 62100 49890 62156
rect 49754 62020 49810 62076
rect 49834 62020 49890 62076
rect 49754 61940 49810 61996
rect 49834 61940 49890 61996
rect 53048 62180 53104 62236
rect 53048 62100 53104 62156
rect 53048 62020 53104 62076
rect 53048 61940 53104 61996
rect 53206 62180 53262 62236
rect 53206 62100 53262 62156
rect 53206 62020 53262 62076
rect 53206 61940 53262 61996
rect 53562 62180 53618 62236
rect 53562 62100 53618 62156
rect 53562 62020 53618 62076
rect 53562 61940 53618 61996
rect 54880 62180 54936 62236
rect 54880 62100 54936 62156
rect 54880 62020 54936 62076
rect 54880 61940 54936 61996
rect 55473 62180 55529 62236
rect 55473 62100 55529 62156
rect 55473 62020 55529 62076
rect 55473 61940 55529 61996
rect 56619 62180 56675 62236
rect 56619 62100 56675 62156
rect 56619 62020 56675 62076
rect 56619 61940 56675 61996
rect 58055 62180 58111 62236
rect 58135 62180 58191 62236
rect 58055 62100 58111 62156
rect 58135 62100 58191 62156
rect 58055 62020 58111 62076
rect 58135 62020 58191 62076
rect 58055 61940 58111 61996
rect 58135 61940 58191 61996
rect 59298 62180 59354 62236
rect 59298 62100 59354 62156
rect 59298 62020 59354 62076
rect 59298 61940 59354 61996
rect 59456 62180 59512 62236
rect 59456 62100 59512 62156
rect 59456 62020 59512 62076
rect 59456 61940 59512 61996
rect 59764 62180 59820 62236
rect 59764 62100 59820 62156
rect 59764 62020 59820 62076
rect 59764 61940 59820 61996
rect 59910 62180 59966 62236
rect 59910 62100 59966 62156
rect 59910 62020 59966 62076
rect 59910 61940 59966 61996
rect 60046 62180 60102 62236
rect 60126 62180 60182 62236
rect 60046 62100 60102 62156
rect 60126 62100 60182 62156
rect 60046 62020 60102 62076
rect 60126 62020 60182 62076
rect 60046 61940 60102 61996
rect 60126 61940 60182 61996
rect 62418 62180 62474 62236
rect 62498 62180 62554 62236
rect 62418 62100 62474 62156
rect 62498 62100 62554 62156
rect 62418 62020 62474 62076
rect 62498 62020 62554 62076
rect 62418 61940 62474 61996
rect 62498 61940 62554 61996
rect 63498 61004 63500 61024
rect 63500 61004 63552 61024
rect 63552 61004 63554 61024
rect 63498 60968 63554 61004
rect 63498 58692 63500 58712
rect 63500 58692 63552 58712
rect 63552 58692 63554 58712
rect 63498 58656 63554 58692
rect 63498 56652 63500 56672
rect 63500 56652 63552 56672
rect 63552 56652 63554 56672
rect 63498 56616 63554 56652
rect 63498 54712 63554 54768
rect 2136 54532 2192 54588
rect 2136 54452 2192 54508
rect 2136 54372 2192 54428
rect 2136 54292 2192 54348
rect 5632 54532 5688 54588
rect 5632 54452 5688 54508
rect 5632 54372 5688 54428
rect 5632 54292 5688 54348
rect 8522 54532 8578 54588
rect 8522 54452 8578 54508
rect 8522 54372 8578 54428
rect 8522 54292 8578 54348
rect 11412 54532 11468 54588
rect 11412 54452 11468 54508
rect 11412 54372 11468 54428
rect 11412 54292 11468 54348
rect 14302 54532 14358 54588
rect 14302 54452 14358 54508
rect 14302 54372 14358 54428
rect 14302 54292 14358 54348
rect 17192 54532 17248 54588
rect 17192 54452 17248 54508
rect 17192 54372 17248 54428
rect 17192 54292 17248 54348
rect 20082 54532 20138 54588
rect 20082 54452 20138 54508
rect 20082 54372 20138 54428
rect 20082 54292 20138 54348
rect 22972 54532 23028 54588
rect 22972 54452 23028 54508
rect 22972 54372 23028 54428
rect 22972 54292 23028 54348
rect 25862 54532 25918 54588
rect 25862 54452 25918 54508
rect 25862 54372 25918 54428
rect 25862 54292 25918 54348
rect 28752 54532 28808 54588
rect 28752 54452 28808 54508
rect 28752 54372 28808 54428
rect 28752 54292 28808 54348
rect 31642 54532 31698 54588
rect 31642 54452 31698 54508
rect 31642 54372 31698 54428
rect 31642 54292 31698 54348
rect 34532 54532 34588 54588
rect 34532 54452 34588 54508
rect 34532 54372 34588 54428
rect 34532 54292 34588 54348
rect 37422 54532 37478 54588
rect 37422 54452 37478 54508
rect 37422 54372 37478 54428
rect 37422 54292 37478 54348
rect 40312 54532 40368 54588
rect 40312 54452 40368 54508
rect 40312 54372 40368 54428
rect 40312 54292 40368 54348
rect 43202 54532 43258 54588
rect 43202 54452 43258 54508
rect 43202 54372 43258 54428
rect 43202 54292 43258 54348
rect 46092 54532 46148 54588
rect 46092 54452 46148 54508
rect 46092 54372 46148 54428
rect 46092 54292 46148 54348
rect 49100 54532 49156 54588
rect 49100 54452 49156 54508
rect 49100 54372 49156 54428
rect 49100 54292 49156 54348
rect 52329 54532 52385 54588
rect 52329 54452 52385 54508
rect 52329 54372 52385 54428
rect 52329 54292 52385 54348
rect 53730 54532 53786 54588
rect 53730 54452 53786 54508
rect 53730 54372 53786 54428
rect 53730 54292 53786 54348
rect 53898 54532 53954 54588
rect 53898 54452 53954 54508
rect 53898 54372 53954 54428
rect 53898 54292 53954 54348
rect 54642 54532 54698 54588
rect 54642 54452 54698 54508
rect 54642 54372 54698 54428
rect 54642 54292 54698 54348
rect 55032 54532 55088 54588
rect 55032 54452 55088 54508
rect 55032 54372 55088 54428
rect 55032 54292 55088 54348
rect 55748 54532 55804 54588
rect 55748 54452 55804 54508
rect 55748 54372 55804 54428
rect 55748 54292 55804 54348
rect 56326 54532 56382 54588
rect 56326 54452 56382 54508
rect 56326 54372 56382 54428
rect 56326 54292 56382 54348
rect 56771 54532 56827 54588
rect 56771 54452 56827 54508
rect 56771 54372 56827 54428
rect 56771 54292 56827 54348
rect 57075 54532 57131 54588
rect 57075 54452 57131 54508
rect 57075 54372 57131 54428
rect 57075 54292 57131 54348
rect 57917 54532 57973 54588
rect 57917 54452 57973 54508
rect 57917 54372 57973 54428
rect 57917 54292 57973 54348
rect 58557 54532 58613 54588
rect 58557 54452 58613 54508
rect 58557 54372 58613 54428
rect 58557 54292 58613 54348
rect 59140 54532 59196 54588
rect 59140 54452 59196 54508
rect 59140 54372 59196 54428
rect 59140 54292 59196 54348
rect 60418 54532 60474 54588
rect 60418 54452 60474 54508
rect 60418 54372 60474 54428
rect 60418 54292 60474 54348
rect 60576 54532 60632 54588
rect 60576 54452 60632 54508
rect 60576 54372 60632 54428
rect 60576 54292 60632 54348
rect 62620 54532 62676 54588
rect 62700 54532 62756 54588
rect 62620 54452 62676 54508
rect 62700 54452 62756 54508
rect 62620 54372 62676 54428
rect 62700 54372 62756 54428
rect 62620 54292 62676 54348
rect 62700 54292 62756 54348
rect 2276 52180 2332 52236
rect 2356 52180 2412 52236
rect 2276 52100 2332 52156
rect 2356 52100 2412 52156
rect 2276 52020 2332 52076
rect 2356 52020 2412 52076
rect 2276 51940 2332 51996
rect 2356 51940 2412 51996
rect 5485 52180 5541 52236
rect 5485 52100 5541 52156
rect 5485 52020 5541 52076
rect 5485 51940 5541 51996
rect 8375 52180 8431 52236
rect 8375 52100 8431 52156
rect 8375 52020 8431 52076
rect 8375 51940 8431 51996
rect 11265 52180 11321 52236
rect 11265 52100 11321 52156
rect 11265 52020 11321 52076
rect 11265 51940 11321 51996
rect 14155 52180 14211 52236
rect 14155 52100 14211 52156
rect 14155 52020 14211 52076
rect 14155 51940 14211 51996
rect 17045 52180 17101 52236
rect 17045 52100 17101 52156
rect 17045 52020 17101 52076
rect 17045 51940 17101 51996
rect 19935 52180 19991 52236
rect 19935 52100 19991 52156
rect 19935 52020 19991 52076
rect 19935 51940 19991 51996
rect 22825 52180 22881 52236
rect 22825 52100 22881 52156
rect 22825 52020 22881 52076
rect 22825 51940 22881 51996
rect 25715 52180 25771 52236
rect 25715 52100 25771 52156
rect 25715 52020 25771 52076
rect 25715 51940 25771 51996
rect 28605 52180 28661 52236
rect 28605 52100 28661 52156
rect 28605 52020 28661 52076
rect 28605 51940 28661 51996
rect 31495 52180 31551 52236
rect 31495 52100 31551 52156
rect 31495 52020 31551 52076
rect 31495 51940 31551 51996
rect 34385 52180 34441 52236
rect 34385 52100 34441 52156
rect 34385 52020 34441 52076
rect 34385 51940 34441 51996
rect 37275 52180 37331 52236
rect 37275 52100 37331 52156
rect 37275 52020 37331 52076
rect 37275 51940 37331 51996
rect 40165 52180 40221 52236
rect 40165 52100 40221 52156
rect 40165 52020 40221 52076
rect 40165 51940 40221 51996
rect 43055 52180 43111 52236
rect 43055 52100 43111 52156
rect 43055 52020 43111 52076
rect 43055 51940 43111 51996
rect 45945 52180 46001 52236
rect 45945 52100 46001 52156
rect 45945 52020 46001 52076
rect 45945 51940 46001 51996
rect 48892 52180 48948 52236
rect 48892 52100 48948 52156
rect 48892 52020 48948 52076
rect 48892 51940 48948 51996
rect 49754 52180 49810 52236
rect 49834 52180 49890 52236
rect 49754 52100 49810 52156
rect 49834 52100 49890 52156
rect 49754 52020 49810 52076
rect 49834 52020 49890 52076
rect 49754 51940 49810 51996
rect 49834 51940 49890 51996
rect 53048 52180 53104 52236
rect 53048 52100 53104 52156
rect 53048 52020 53104 52076
rect 53048 51940 53104 51996
rect 53206 52180 53262 52236
rect 53206 52100 53262 52156
rect 53206 52020 53262 52076
rect 53206 51940 53262 51996
rect 53562 52180 53618 52236
rect 53562 52100 53618 52156
rect 53562 52020 53618 52076
rect 53562 51940 53618 51996
rect 54880 52180 54936 52236
rect 54880 52100 54936 52156
rect 54880 52020 54936 52076
rect 54880 51940 54936 51996
rect 55473 52180 55529 52236
rect 55473 52100 55529 52156
rect 55473 52020 55529 52076
rect 55473 51940 55529 51996
rect 56619 52180 56675 52236
rect 56619 52100 56675 52156
rect 56619 52020 56675 52076
rect 56619 51940 56675 51996
rect 58055 52180 58111 52236
rect 58135 52180 58191 52236
rect 58055 52100 58111 52156
rect 58135 52100 58191 52156
rect 58055 52020 58111 52076
rect 58135 52020 58191 52076
rect 58055 51940 58111 51996
rect 58135 51940 58191 51996
rect 59298 52180 59354 52236
rect 59298 52100 59354 52156
rect 59298 52020 59354 52076
rect 59298 51940 59354 51996
rect 59456 52180 59512 52236
rect 59456 52100 59512 52156
rect 59456 52020 59512 52076
rect 59456 51940 59512 51996
rect 59764 52180 59820 52236
rect 59764 52100 59820 52156
rect 59764 52020 59820 52076
rect 59764 51940 59820 51996
rect 59910 52180 59966 52236
rect 59910 52100 59966 52156
rect 59910 52020 59966 52076
rect 59910 51940 59966 51996
rect 60046 52180 60102 52236
rect 60126 52180 60182 52236
rect 60046 52100 60102 52156
rect 60126 52100 60182 52156
rect 60046 52020 60102 52076
rect 60126 52020 60182 52076
rect 60046 51940 60102 51996
rect 60126 51940 60182 51996
rect 62418 52180 62474 52236
rect 62498 52180 62554 52236
rect 62418 52100 62474 52156
rect 62498 52100 62554 52156
rect 62418 52020 62474 52076
rect 62498 52020 62554 52076
rect 62418 51940 62474 51996
rect 62498 51940 62554 51996
rect 2136 44532 2192 44588
rect 2136 44452 2192 44508
rect 2136 44372 2192 44428
rect 2136 44292 2192 44348
rect 5632 44532 5688 44588
rect 5632 44452 5688 44508
rect 5632 44372 5688 44428
rect 5632 44292 5688 44348
rect 8522 44532 8578 44588
rect 8522 44452 8578 44508
rect 8522 44372 8578 44428
rect 8522 44292 8578 44348
rect 11412 44532 11468 44588
rect 11412 44452 11468 44508
rect 11412 44372 11468 44428
rect 11412 44292 11468 44348
rect 14302 44532 14358 44588
rect 14302 44452 14358 44508
rect 14302 44372 14358 44428
rect 14302 44292 14358 44348
rect 17192 44532 17248 44588
rect 17192 44452 17248 44508
rect 17192 44372 17248 44428
rect 17192 44292 17248 44348
rect 20082 44532 20138 44588
rect 20082 44452 20138 44508
rect 20082 44372 20138 44428
rect 20082 44292 20138 44348
rect 22972 44532 23028 44588
rect 22972 44452 23028 44508
rect 22972 44372 23028 44428
rect 22972 44292 23028 44348
rect 25862 44532 25918 44588
rect 25862 44452 25918 44508
rect 25862 44372 25918 44428
rect 25862 44292 25918 44348
rect 28752 44532 28808 44588
rect 28752 44452 28808 44508
rect 28752 44372 28808 44428
rect 28752 44292 28808 44348
rect 31642 44532 31698 44588
rect 31642 44452 31698 44508
rect 31642 44372 31698 44428
rect 31642 44292 31698 44348
rect 34532 44532 34588 44588
rect 34532 44452 34588 44508
rect 34532 44372 34588 44428
rect 34532 44292 34588 44348
rect 37422 44532 37478 44588
rect 37422 44452 37478 44508
rect 37422 44372 37478 44428
rect 37422 44292 37478 44348
rect 40312 44532 40368 44588
rect 40312 44452 40368 44508
rect 40312 44372 40368 44428
rect 40312 44292 40368 44348
rect 43202 44532 43258 44588
rect 43202 44452 43258 44508
rect 43202 44372 43258 44428
rect 43202 44292 43258 44348
rect 46092 44532 46148 44588
rect 46092 44452 46148 44508
rect 46092 44372 46148 44428
rect 46092 44292 46148 44348
rect 52329 44532 52385 44588
rect 52329 44452 52385 44508
rect 52329 44372 52385 44428
rect 52329 44292 52385 44348
rect 53730 44532 53786 44588
rect 53730 44452 53786 44508
rect 53730 44372 53786 44428
rect 53730 44292 53786 44348
rect 54642 44532 54698 44588
rect 54642 44452 54698 44508
rect 54642 44372 54698 44428
rect 54642 44292 54698 44348
rect 55032 44532 55088 44588
rect 55032 44452 55088 44508
rect 55032 44372 55088 44428
rect 55032 44292 55088 44348
rect 55748 44532 55804 44588
rect 55748 44452 55804 44508
rect 55748 44372 55804 44428
rect 55748 44292 55804 44348
rect 56326 44532 56382 44588
rect 56326 44452 56382 44508
rect 56326 44372 56382 44428
rect 56326 44292 56382 44348
rect 56771 44532 56827 44588
rect 56771 44452 56827 44508
rect 56771 44372 56827 44428
rect 56771 44292 56827 44348
rect 57075 44532 57131 44588
rect 57075 44452 57131 44508
rect 57075 44372 57131 44428
rect 57075 44292 57131 44348
rect 57917 44532 57973 44588
rect 57917 44452 57973 44508
rect 57917 44372 57973 44428
rect 57917 44292 57973 44348
rect 58441 44532 58497 44588
rect 58441 44452 58497 44508
rect 58441 44372 58497 44428
rect 58441 44292 58497 44348
rect 59140 44532 59196 44588
rect 59140 44452 59196 44508
rect 59140 44372 59196 44428
rect 59140 44292 59196 44348
rect 60418 44532 60474 44588
rect 60418 44452 60474 44508
rect 60418 44372 60474 44428
rect 60418 44292 60474 44348
rect 60576 44532 60632 44588
rect 60576 44452 60632 44508
rect 60576 44372 60632 44428
rect 60576 44292 60632 44348
rect 62620 44532 62676 44588
rect 62700 44532 62756 44588
rect 62620 44452 62676 44508
rect 62700 44452 62756 44508
rect 62620 44372 62676 44428
rect 62700 44372 62756 44428
rect 62620 44292 62676 44348
rect 62700 44292 62756 44348
rect 2276 42180 2332 42236
rect 2356 42180 2412 42236
rect 2276 42100 2332 42156
rect 2356 42100 2412 42156
rect 2276 42020 2332 42076
rect 2356 42020 2412 42076
rect 2276 41940 2332 41996
rect 2356 41940 2412 41996
rect 5485 42180 5541 42236
rect 5485 42100 5541 42156
rect 5485 42020 5541 42076
rect 5485 41940 5541 41996
rect 8375 42180 8431 42236
rect 8375 42100 8431 42156
rect 8375 42020 8431 42076
rect 8375 41940 8431 41996
rect 11265 42180 11321 42236
rect 11265 42100 11321 42156
rect 11265 42020 11321 42076
rect 11265 41940 11321 41996
rect 14155 42180 14211 42236
rect 14155 42100 14211 42156
rect 14155 42020 14211 42076
rect 14155 41940 14211 41996
rect 17045 42180 17101 42236
rect 17045 42100 17101 42156
rect 17045 42020 17101 42076
rect 17045 41940 17101 41996
rect 19935 42180 19991 42236
rect 19935 42100 19991 42156
rect 19935 42020 19991 42076
rect 19935 41940 19991 41996
rect 22825 42180 22881 42236
rect 22825 42100 22881 42156
rect 22825 42020 22881 42076
rect 22825 41940 22881 41996
rect 25715 42180 25771 42236
rect 25715 42100 25771 42156
rect 25715 42020 25771 42076
rect 25715 41940 25771 41996
rect 28605 42180 28661 42236
rect 28605 42100 28661 42156
rect 28605 42020 28661 42076
rect 28605 41940 28661 41996
rect 31495 42180 31551 42236
rect 31495 42100 31551 42156
rect 31495 42020 31551 42076
rect 31495 41940 31551 41996
rect 34385 42180 34441 42236
rect 34385 42100 34441 42156
rect 34385 42020 34441 42076
rect 34385 41940 34441 41996
rect 37275 42180 37331 42236
rect 37275 42100 37331 42156
rect 37275 42020 37331 42076
rect 37275 41940 37331 41996
rect 40165 42180 40221 42236
rect 40165 42100 40221 42156
rect 40165 42020 40221 42076
rect 40165 41940 40221 41996
rect 43055 42180 43111 42236
rect 43055 42100 43111 42156
rect 43055 42020 43111 42076
rect 43055 41940 43111 41996
rect 45945 42180 46001 42236
rect 45945 42100 46001 42156
rect 45945 42020 46001 42076
rect 45945 41940 46001 41996
rect 48892 42180 48948 42236
rect 48892 42100 48948 42156
rect 48892 42020 48948 42076
rect 48892 41940 48948 41996
rect 49754 42180 49810 42236
rect 49834 42180 49890 42236
rect 49754 42100 49810 42156
rect 49834 42100 49890 42156
rect 49754 42020 49810 42076
rect 49834 42020 49890 42076
rect 49754 41940 49810 41996
rect 49834 41940 49890 41996
rect 53048 42180 53104 42236
rect 53048 42100 53104 42156
rect 53048 42020 53104 42076
rect 53048 41940 53104 41996
rect 53206 42180 53262 42236
rect 53206 42100 53262 42156
rect 53206 42020 53262 42076
rect 53206 41940 53262 41996
rect 53562 42180 53618 42236
rect 53562 42100 53618 42156
rect 53562 42020 53618 42076
rect 53562 41940 53618 41996
rect 54880 42180 54936 42236
rect 54880 42100 54936 42156
rect 54880 42020 54936 42076
rect 54880 41940 54936 41996
rect 55473 42180 55529 42236
rect 55473 42100 55529 42156
rect 55473 42020 55529 42076
rect 55473 41940 55529 41996
rect 56619 42180 56675 42236
rect 56619 42100 56675 42156
rect 56619 42020 56675 42076
rect 56619 41940 56675 41996
rect 58055 42180 58111 42236
rect 58135 42180 58191 42236
rect 58055 42100 58111 42156
rect 58135 42100 58191 42156
rect 58055 42020 58111 42076
rect 58135 42020 58191 42076
rect 58055 41940 58111 41996
rect 58135 41940 58191 41996
rect 59298 42180 59354 42236
rect 59298 42100 59354 42156
rect 59298 42020 59354 42076
rect 59298 41940 59354 41996
rect 59456 42180 59512 42236
rect 59456 42100 59512 42156
rect 59456 42020 59512 42076
rect 59456 41940 59512 41996
rect 59764 42180 59820 42236
rect 59764 42100 59820 42156
rect 59764 42020 59820 42076
rect 59764 41940 59820 41996
rect 59910 42180 59966 42236
rect 59910 42100 59966 42156
rect 59910 42020 59966 42076
rect 59910 41940 59966 41996
rect 60046 42180 60102 42236
rect 60126 42180 60182 42236
rect 60046 42100 60102 42156
rect 60126 42100 60182 42156
rect 60046 42020 60102 42076
rect 60126 42020 60182 42076
rect 60046 41940 60102 41996
rect 60126 41940 60182 41996
rect 62418 42180 62474 42236
rect 62498 42180 62554 42236
rect 62418 42100 62474 42156
rect 62498 42100 62554 42156
rect 62418 42020 62474 42076
rect 62498 42020 62554 42076
rect 62418 41940 62474 41996
rect 62498 41940 62554 41996
rect 2136 34532 2192 34588
rect 2136 34452 2192 34508
rect 2136 34372 2192 34428
rect 2136 34292 2192 34348
rect 5632 34532 5688 34588
rect 5632 34452 5688 34508
rect 5632 34372 5688 34428
rect 5632 34292 5688 34348
rect 8522 34532 8578 34588
rect 8522 34452 8578 34508
rect 8522 34372 8578 34428
rect 8522 34292 8578 34348
rect 11412 34532 11468 34588
rect 11412 34452 11468 34508
rect 11412 34372 11468 34428
rect 11412 34292 11468 34348
rect 14302 34532 14358 34588
rect 14302 34452 14358 34508
rect 14302 34372 14358 34428
rect 14302 34292 14358 34348
rect 17192 34532 17248 34588
rect 17192 34452 17248 34508
rect 17192 34372 17248 34428
rect 17192 34292 17248 34348
rect 20082 34532 20138 34588
rect 20082 34452 20138 34508
rect 20082 34372 20138 34428
rect 20082 34292 20138 34348
rect 22972 34532 23028 34588
rect 22972 34452 23028 34508
rect 22972 34372 23028 34428
rect 22972 34292 23028 34348
rect 25862 34532 25918 34588
rect 25862 34452 25918 34508
rect 25862 34372 25918 34428
rect 25862 34292 25918 34348
rect 28752 34532 28808 34588
rect 28752 34452 28808 34508
rect 28752 34372 28808 34428
rect 28752 34292 28808 34348
rect 31642 34532 31698 34588
rect 31642 34452 31698 34508
rect 31642 34372 31698 34428
rect 31642 34292 31698 34348
rect 34532 34532 34588 34588
rect 34532 34452 34588 34508
rect 34532 34372 34588 34428
rect 34532 34292 34588 34348
rect 37422 34532 37478 34588
rect 37422 34452 37478 34508
rect 37422 34372 37478 34428
rect 37422 34292 37478 34348
rect 40312 34532 40368 34588
rect 40312 34452 40368 34508
rect 40312 34372 40368 34428
rect 40312 34292 40368 34348
rect 43202 34532 43258 34588
rect 43202 34452 43258 34508
rect 43202 34372 43258 34428
rect 43202 34292 43258 34348
rect 46092 34532 46148 34588
rect 46092 34452 46148 34508
rect 46092 34372 46148 34428
rect 46092 34292 46148 34348
rect 49100 34532 49156 34588
rect 49100 34452 49156 34508
rect 49100 34372 49156 34428
rect 49100 34292 49156 34348
rect 52329 34532 52385 34588
rect 52329 34452 52385 34508
rect 52329 34372 52385 34428
rect 52329 34292 52385 34348
rect 53730 34532 53786 34588
rect 53730 34452 53786 34508
rect 53730 34372 53786 34428
rect 53730 34292 53786 34348
rect 53898 34532 53954 34588
rect 53898 34452 53954 34508
rect 53898 34372 53954 34428
rect 53898 34292 53954 34348
rect 54642 34532 54698 34588
rect 54642 34452 54698 34508
rect 54642 34372 54698 34428
rect 54642 34292 54698 34348
rect 55032 34532 55088 34588
rect 55032 34452 55088 34508
rect 55032 34372 55088 34428
rect 55032 34292 55088 34348
rect 55748 34532 55804 34588
rect 55748 34452 55804 34508
rect 55748 34372 55804 34428
rect 55748 34292 55804 34348
rect 56326 34532 56382 34588
rect 56326 34452 56382 34508
rect 56326 34372 56382 34428
rect 56326 34292 56382 34348
rect 56771 34532 56827 34588
rect 56771 34452 56827 34508
rect 56771 34372 56827 34428
rect 56771 34292 56827 34348
rect 57075 34532 57131 34588
rect 57075 34452 57131 34508
rect 57075 34372 57131 34428
rect 57075 34292 57131 34348
rect 57917 34532 57973 34588
rect 57917 34452 57973 34508
rect 57917 34372 57973 34428
rect 57917 34292 57973 34348
rect 58557 34532 58613 34588
rect 58557 34452 58613 34508
rect 58557 34372 58613 34428
rect 58557 34292 58613 34348
rect 59140 34532 59196 34588
rect 59140 34452 59196 34508
rect 59140 34372 59196 34428
rect 59140 34292 59196 34348
rect 60418 34532 60474 34588
rect 60418 34452 60474 34508
rect 60418 34372 60474 34428
rect 60418 34292 60474 34348
rect 60576 34532 60632 34588
rect 60576 34452 60632 34508
rect 60576 34372 60632 34428
rect 60576 34292 60632 34348
rect 62620 34532 62676 34588
rect 62700 34532 62756 34588
rect 62620 34452 62676 34508
rect 62700 34452 62756 34508
rect 62620 34372 62676 34428
rect 62700 34372 62756 34428
rect 62620 34292 62676 34348
rect 62700 34292 62756 34348
rect 2276 32180 2332 32236
rect 2356 32180 2412 32236
rect 2276 32100 2332 32156
rect 2356 32100 2412 32156
rect 2276 32020 2332 32076
rect 2356 32020 2412 32076
rect 2276 31940 2332 31996
rect 2356 31940 2412 31996
rect 5485 32180 5541 32236
rect 5485 32100 5541 32156
rect 5485 32020 5541 32076
rect 5485 31940 5541 31996
rect 8375 32180 8431 32236
rect 8375 32100 8431 32156
rect 8375 32020 8431 32076
rect 8375 31940 8431 31996
rect 11265 32180 11321 32236
rect 11265 32100 11321 32156
rect 11265 32020 11321 32076
rect 11265 31940 11321 31996
rect 14155 32180 14211 32236
rect 14155 32100 14211 32156
rect 14155 32020 14211 32076
rect 14155 31940 14211 31996
rect 17045 32180 17101 32236
rect 17045 32100 17101 32156
rect 17045 32020 17101 32076
rect 17045 31940 17101 31996
rect 19935 32180 19991 32236
rect 19935 32100 19991 32156
rect 19935 32020 19991 32076
rect 19935 31940 19991 31996
rect 22825 32180 22881 32236
rect 22825 32100 22881 32156
rect 22825 32020 22881 32076
rect 22825 31940 22881 31996
rect 25715 32180 25771 32236
rect 25715 32100 25771 32156
rect 25715 32020 25771 32076
rect 25715 31940 25771 31996
rect 28605 32180 28661 32236
rect 28605 32100 28661 32156
rect 28605 32020 28661 32076
rect 28605 31940 28661 31996
rect 31495 32180 31551 32236
rect 31495 32100 31551 32156
rect 31495 32020 31551 32076
rect 31495 31940 31551 31996
rect 34385 32180 34441 32236
rect 34385 32100 34441 32156
rect 34385 32020 34441 32076
rect 34385 31940 34441 31996
rect 37275 32180 37331 32236
rect 37275 32100 37331 32156
rect 37275 32020 37331 32076
rect 37275 31940 37331 31996
rect 40165 32180 40221 32236
rect 40165 32100 40221 32156
rect 40165 32020 40221 32076
rect 40165 31940 40221 31996
rect 43055 32180 43111 32236
rect 43055 32100 43111 32156
rect 43055 32020 43111 32076
rect 43055 31940 43111 31996
rect 45945 32180 46001 32236
rect 45945 32100 46001 32156
rect 45945 32020 46001 32076
rect 45945 31940 46001 31996
rect 48892 32180 48948 32236
rect 48892 32100 48948 32156
rect 48892 32020 48948 32076
rect 48892 31940 48948 31996
rect 49754 32180 49810 32236
rect 49834 32180 49890 32236
rect 49754 32100 49810 32156
rect 49834 32100 49890 32156
rect 49754 32020 49810 32076
rect 49834 32020 49890 32076
rect 49754 31940 49810 31996
rect 49834 31940 49890 31996
rect 53048 32180 53104 32236
rect 53048 32100 53104 32156
rect 53048 32020 53104 32076
rect 53048 31940 53104 31996
rect 53206 32180 53262 32236
rect 53206 32100 53262 32156
rect 53206 32020 53262 32076
rect 53206 31940 53262 31996
rect 53562 32180 53618 32236
rect 53562 32100 53618 32156
rect 53562 32020 53618 32076
rect 53562 31940 53618 31996
rect 54880 32180 54936 32236
rect 54880 32100 54936 32156
rect 54880 32020 54936 32076
rect 54880 31940 54936 31996
rect 55473 32180 55529 32236
rect 55473 32100 55529 32156
rect 55473 32020 55529 32076
rect 55473 31940 55529 31996
rect 56619 32180 56675 32236
rect 56619 32100 56675 32156
rect 56619 32020 56675 32076
rect 56619 31940 56675 31996
rect 58055 32180 58111 32236
rect 58135 32180 58191 32236
rect 58055 32100 58111 32156
rect 58135 32100 58191 32156
rect 58055 32020 58111 32076
rect 58135 32020 58191 32076
rect 58055 31940 58111 31996
rect 58135 31940 58191 31996
rect 59298 32180 59354 32236
rect 59298 32100 59354 32156
rect 59298 32020 59354 32076
rect 59298 31940 59354 31996
rect 59456 32180 59512 32236
rect 59456 32100 59512 32156
rect 59456 32020 59512 32076
rect 59456 31940 59512 31996
rect 59764 32180 59820 32236
rect 59764 32100 59820 32156
rect 59764 32020 59820 32076
rect 59764 31940 59820 31996
rect 59910 32180 59966 32236
rect 59910 32100 59966 32156
rect 59910 32020 59966 32076
rect 59910 31940 59966 31996
rect 60046 32180 60102 32236
rect 60126 32180 60182 32236
rect 60046 32100 60102 32156
rect 60126 32100 60182 32156
rect 60046 32020 60102 32076
rect 60126 32020 60182 32076
rect 60046 31940 60102 31996
rect 60126 31940 60182 31996
rect 62418 32180 62474 32236
rect 62498 32180 62554 32236
rect 62418 32100 62474 32156
rect 62498 32100 62554 32156
rect 62418 32020 62474 32076
rect 62498 32020 62554 32076
rect 62418 31940 62474 31996
rect 62498 31940 62554 31996
rect 2136 24532 2192 24588
rect 2136 24452 2192 24508
rect 2136 24372 2192 24428
rect 2136 24292 2192 24348
rect 5632 24532 5688 24588
rect 5632 24452 5688 24508
rect 5632 24372 5688 24428
rect 5632 24292 5688 24348
rect 8522 24532 8578 24588
rect 8522 24452 8578 24508
rect 8522 24372 8578 24428
rect 8522 24292 8578 24348
rect 11412 24532 11468 24588
rect 11412 24452 11468 24508
rect 11412 24372 11468 24428
rect 11412 24292 11468 24348
rect 14302 24532 14358 24588
rect 14302 24452 14358 24508
rect 14302 24372 14358 24428
rect 14302 24292 14358 24348
rect 17192 24532 17248 24588
rect 17192 24452 17248 24508
rect 17192 24372 17248 24428
rect 17192 24292 17248 24348
rect 20082 24532 20138 24588
rect 20082 24452 20138 24508
rect 20082 24372 20138 24428
rect 20082 24292 20138 24348
rect 22972 24532 23028 24588
rect 22972 24452 23028 24508
rect 22972 24372 23028 24428
rect 22972 24292 23028 24348
rect 25862 24532 25918 24588
rect 25862 24452 25918 24508
rect 25862 24372 25918 24428
rect 25862 24292 25918 24348
rect 28752 24532 28808 24588
rect 28752 24452 28808 24508
rect 28752 24372 28808 24428
rect 28752 24292 28808 24348
rect 31642 24532 31698 24588
rect 31642 24452 31698 24508
rect 31642 24372 31698 24428
rect 31642 24292 31698 24348
rect 34532 24532 34588 24588
rect 34532 24452 34588 24508
rect 34532 24372 34588 24428
rect 34532 24292 34588 24348
rect 37422 24532 37478 24588
rect 37422 24452 37478 24508
rect 37422 24372 37478 24428
rect 37422 24292 37478 24348
rect 40312 24532 40368 24588
rect 40312 24452 40368 24508
rect 40312 24372 40368 24428
rect 40312 24292 40368 24348
rect 43202 24532 43258 24588
rect 43202 24452 43258 24508
rect 43202 24372 43258 24428
rect 43202 24292 43258 24348
rect 46092 24532 46148 24588
rect 46092 24452 46148 24508
rect 46092 24372 46148 24428
rect 46092 24292 46148 24348
rect 49100 24532 49156 24588
rect 49100 24452 49156 24508
rect 49100 24372 49156 24428
rect 49100 24292 49156 24348
rect 52329 24532 52385 24588
rect 52329 24452 52385 24508
rect 52329 24372 52385 24428
rect 52329 24292 52385 24348
rect 53730 24532 53786 24588
rect 53730 24452 53786 24508
rect 53730 24372 53786 24428
rect 53730 24292 53786 24348
rect 53898 24532 53954 24588
rect 53898 24452 53954 24508
rect 53898 24372 53954 24428
rect 53898 24292 53954 24348
rect 54642 24532 54698 24588
rect 54642 24452 54698 24508
rect 54642 24372 54698 24428
rect 54642 24292 54698 24348
rect 55032 24532 55088 24588
rect 55032 24452 55088 24508
rect 55032 24372 55088 24428
rect 55032 24292 55088 24348
rect 55748 24532 55804 24588
rect 55748 24452 55804 24508
rect 55748 24372 55804 24428
rect 55748 24292 55804 24348
rect 56326 24532 56382 24588
rect 56326 24452 56382 24508
rect 56326 24372 56382 24428
rect 56326 24292 56382 24348
rect 56771 24532 56827 24588
rect 56771 24452 56827 24508
rect 56771 24372 56827 24428
rect 56771 24292 56827 24348
rect 57075 24532 57131 24588
rect 57075 24452 57131 24508
rect 57075 24372 57131 24428
rect 57075 24292 57131 24348
rect 57917 24532 57973 24588
rect 57917 24452 57973 24508
rect 57917 24372 57973 24428
rect 57917 24292 57973 24348
rect 58557 24532 58613 24588
rect 58557 24452 58613 24508
rect 58557 24372 58613 24428
rect 58557 24292 58613 24348
rect 59140 24532 59196 24588
rect 59140 24452 59196 24508
rect 59140 24372 59196 24428
rect 59140 24292 59196 24348
rect 60418 24532 60474 24588
rect 60418 24452 60474 24508
rect 60418 24372 60474 24428
rect 60418 24292 60474 24348
rect 60576 24532 60632 24588
rect 60576 24452 60632 24508
rect 60576 24372 60632 24428
rect 60576 24292 60632 24348
rect 62620 24532 62676 24588
rect 62700 24532 62756 24588
rect 62620 24452 62676 24508
rect 62700 24452 62756 24508
rect 62620 24372 62676 24428
rect 62700 24372 62756 24428
rect 62620 24292 62676 24348
rect 62700 24292 62756 24348
rect 2276 22180 2332 22236
rect 2356 22180 2412 22236
rect 2276 22100 2332 22156
rect 2356 22100 2412 22156
rect 2276 22020 2332 22076
rect 2356 22020 2412 22076
rect 2276 21940 2332 21996
rect 2356 21940 2412 21996
rect 5485 22180 5541 22236
rect 5485 22100 5541 22156
rect 5485 22020 5541 22076
rect 5485 21940 5541 21996
rect 8375 22180 8431 22236
rect 8375 22100 8431 22156
rect 8375 22020 8431 22076
rect 8375 21940 8431 21996
rect 11265 22180 11321 22236
rect 11265 22100 11321 22156
rect 11265 22020 11321 22076
rect 11265 21940 11321 21996
rect 14155 22180 14211 22236
rect 14155 22100 14211 22156
rect 14155 22020 14211 22076
rect 14155 21940 14211 21996
rect 17045 22180 17101 22236
rect 17045 22100 17101 22156
rect 17045 22020 17101 22076
rect 17045 21940 17101 21996
rect 19935 22180 19991 22236
rect 19935 22100 19991 22156
rect 19935 22020 19991 22076
rect 19935 21940 19991 21996
rect 22825 22180 22881 22236
rect 22825 22100 22881 22156
rect 22825 22020 22881 22076
rect 22825 21940 22881 21996
rect 25715 22180 25771 22236
rect 25715 22100 25771 22156
rect 25715 22020 25771 22076
rect 25715 21940 25771 21996
rect 28605 22180 28661 22236
rect 28605 22100 28661 22156
rect 28605 22020 28661 22076
rect 28605 21940 28661 21996
rect 31495 22180 31551 22236
rect 31495 22100 31551 22156
rect 31495 22020 31551 22076
rect 31495 21940 31551 21996
rect 34385 22180 34441 22236
rect 34385 22100 34441 22156
rect 34385 22020 34441 22076
rect 34385 21940 34441 21996
rect 37275 22180 37331 22236
rect 37275 22100 37331 22156
rect 37275 22020 37331 22076
rect 37275 21940 37331 21996
rect 40165 22180 40221 22236
rect 40165 22100 40221 22156
rect 40165 22020 40221 22076
rect 40165 21940 40221 21996
rect 43055 22180 43111 22236
rect 43055 22100 43111 22156
rect 43055 22020 43111 22076
rect 43055 21940 43111 21996
rect 45945 22180 46001 22236
rect 45945 22100 46001 22156
rect 45945 22020 46001 22076
rect 45945 21940 46001 21996
rect 48892 22180 48948 22236
rect 48892 22100 48948 22156
rect 48892 22020 48948 22076
rect 48892 21940 48948 21996
rect 49754 22180 49810 22236
rect 49834 22180 49890 22236
rect 49754 22100 49810 22156
rect 49834 22100 49890 22156
rect 49754 22020 49810 22076
rect 49834 22020 49890 22076
rect 49754 21940 49810 21996
rect 49834 21940 49890 21996
rect 53048 22180 53104 22236
rect 53048 22100 53104 22156
rect 53048 22020 53104 22076
rect 53048 21940 53104 21996
rect 53206 22180 53262 22236
rect 53206 22100 53262 22156
rect 53206 22020 53262 22076
rect 53206 21940 53262 21996
rect 53562 22180 53618 22236
rect 53562 22100 53618 22156
rect 53562 22020 53618 22076
rect 53562 21940 53618 21996
rect 54880 22180 54936 22236
rect 54880 22100 54936 22156
rect 54880 22020 54936 22076
rect 54880 21940 54936 21996
rect 55473 22180 55529 22236
rect 55473 22100 55529 22156
rect 55473 22020 55529 22076
rect 55473 21940 55529 21996
rect 56619 22180 56675 22236
rect 56619 22100 56675 22156
rect 56619 22020 56675 22076
rect 56619 21940 56675 21996
rect 58055 22180 58111 22236
rect 58135 22180 58191 22236
rect 58055 22100 58111 22156
rect 58135 22100 58191 22156
rect 58055 22020 58111 22076
rect 58135 22020 58191 22076
rect 58055 21940 58111 21996
rect 58135 21940 58191 21996
rect 59298 22180 59354 22236
rect 59298 22100 59354 22156
rect 59298 22020 59354 22076
rect 59298 21940 59354 21996
rect 59456 22180 59512 22236
rect 59456 22100 59512 22156
rect 59456 22020 59512 22076
rect 59456 21940 59512 21996
rect 59764 22180 59820 22236
rect 59764 22100 59820 22156
rect 59764 22020 59820 22076
rect 59764 21940 59820 21996
rect 59910 22180 59966 22236
rect 59910 22100 59966 22156
rect 59910 22020 59966 22076
rect 59910 21940 59966 21996
rect 60046 22180 60102 22236
rect 60126 22180 60182 22236
rect 60046 22100 60102 22156
rect 60126 22100 60182 22156
rect 60046 22020 60102 22076
rect 60126 22020 60182 22076
rect 60046 21940 60102 21996
rect 60126 21940 60182 21996
rect 62418 22180 62474 22236
rect 62498 22180 62554 22236
rect 62418 22100 62474 22156
rect 62498 22100 62554 22156
rect 62418 22020 62474 22076
rect 62498 22020 62554 22076
rect 62418 21940 62474 21996
rect 62498 21940 62554 21996
rect 2136 14532 2192 14588
rect 2136 14452 2192 14508
rect 2136 14372 2192 14428
rect 2136 14292 2192 14348
rect 5632 14532 5688 14588
rect 5632 14452 5688 14508
rect 5632 14372 5688 14428
rect 5632 14292 5688 14348
rect 8522 14532 8578 14588
rect 8522 14452 8578 14508
rect 8522 14372 8578 14428
rect 8522 14292 8578 14348
rect 11412 14532 11468 14588
rect 11412 14452 11468 14508
rect 11412 14372 11468 14428
rect 11412 14292 11468 14348
rect 14302 14532 14358 14588
rect 14302 14452 14358 14508
rect 14302 14372 14358 14428
rect 14302 14292 14358 14348
rect 17192 14532 17248 14588
rect 17192 14452 17248 14508
rect 17192 14372 17248 14428
rect 17192 14292 17248 14348
rect 20082 14532 20138 14588
rect 20082 14452 20138 14508
rect 20082 14372 20138 14428
rect 20082 14292 20138 14348
rect 22972 14532 23028 14588
rect 22972 14452 23028 14508
rect 22972 14372 23028 14428
rect 22972 14292 23028 14348
rect 25862 14532 25918 14588
rect 25862 14452 25918 14508
rect 25862 14372 25918 14428
rect 25862 14292 25918 14348
rect 28752 14532 28808 14588
rect 28752 14452 28808 14508
rect 28752 14372 28808 14428
rect 28752 14292 28808 14348
rect 31642 14532 31698 14588
rect 31642 14452 31698 14508
rect 31642 14372 31698 14428
rect 31642 14292 31698 14348
rect 34532 14532 34588 14588
rect 34532 14452 34588 14508
rect 34532 14372 34588 14428
rect 34532 14292 34588 14348
rect 37422 14532 37478 14588
rect 37422 14452 37478 14508
rect 37422 14372 37478 14428
rect 37422 14292 37478 14348
rect 40312 14532 40368 14588
rect 40312 14452 40368 14508
rect 40312 14372 40368 14428
rect 40312 14292 40368 14348
rect 43202 14532 43258 14588
rect 43202 14452 43258 14508
rect 43202 14372 43258 14428
rect 43202 14292 43258 14348
rect 46092 14532 46148 14588
rect 46092 14452 46148 14508
rect 46092 14372 46148 14428
rect 46092 14292 46148 14348
rect 49100 14532 49156 14588
rect 49100 14452 49156 14508
rect 49100 14372 49156 14428
rect 49100 14292 49156 14348
rect 52329 14532 52385 14588
rect 52329 14452 52385 14508
rect 52329 14372 52385 14428
rect 52329 14292 52385 14348
rect 53730 14532 53786 14588
rect 53730 14452 53786 14508
rect 53730 14372 53786 14428
rect 53730 14292 53786 14348
rect 53898 14532 53954 14588
rect 53898 14452 53954 14508
rect 53898 14372 53954 14428
rect 53898 14292 53954 14348
rect 54642 14532 54698 14588
rect 54642 14452 54698 14508
rect 54642 14372 54698 14428
rect 54642 14292 54698 14348
rect 55032 14532 55088 14588
rect 55032 14452 55088 14508
rect 55032 14372 55088 14428
rect 55032 14292 55088 14348
rect 55748 14532 55804 14588
rect 55748 14452 55804 14508
rect 55748 14372 55804 14428
rect 55748 14292 55804 14348
rect 56326 14532 56382 14588
rect 56326 14452 56382 14508
rect 56326 14372 56382 14428
rect 56326 14292 56382 14348
rect 56771 14532 56827 14588
rect 56771 14452 56827 14508
rect 56771 14372 56827 14428
rect 56771 14292 56827 14348
rect 57075 14532 57131 14588
rect 57075 14452 57131 14508
rect 57075 14372 57131 14428
rect 57075 14292 57131 14348
rect 57917 14532 57973 14588
rect 57917 14452 57973 14508
rect 57917 14372 57973 14428
rect 57917 14292 57973 14348
rect 58557 14532 58613 14588
rect 58557 14452 58613 14508
rect 58557 14372 58613 14428
rect 58557 14292 58613 14348
rect 59140 14532 59196 14588
rect 59140 14452 59196 14508
rect 59140 14372 59196 14428
rect 59140 14292 59196 14348
rect 60418 14532 60474 14588
rect 60418 14452 60474 14508
rect 60418 14372 60474 14428
rect 60418 14292 60474 14348
rect 60576 14532 60632 14588
rect 60576 14452 60632 14508
rect 60576 14372 60632 14428
rect 60576 14292 60632 14348
rect 62620 14532 62676 14588
rect 62700 14532 62756 14588
rect 62620 14452 62676 14508
rect 62700 14452 62756 14508
rect 62620 14372 62676 14428
rect 62700 14372 62756 14428
rect 62620 14292 62676 14348
rect 62700 14292 62756 14348
rect 2276 12180 2332 12236
rect 2356 12180 2412 12236
rect 2276 12100 2332 12156
rect 2356 12100 2412 12156
rect 2276 12020 2332 12076
rect 2356 12020 2412 12076
rect 2276 11940 2332 11996
rect 2356 11940 2412 11996
rect 5485 12180 5541 12236
rect 5485 12100 5541 12156
rect 5485 12020 5541 12076
rect 5485 11940 5541 11996
rect 8375 12180 8431 12236
rect 8375 12100 8431 12156
rect 8375 12020 8431 12076
rect 8375 11940 8431 11996
rect 11265 12180 11321 12236
rect 11265 12100 11321 12156
rect 11265 12020 11321 12076
rect 11265 11940 11321 11996
rect 14155 12180 14211 12236
rect 14155 12100 14211 12156
rect 14155 12020 14211 12076
rect 14155 11940 14211 11996
rect 17045 12180 17101 12236
rect 17045 12100 17101 12156
rect 17045 12020 17101 12076
rect 17045 11940 17101 11996
rect 19935 12180 19991 12236
rect 19935 12100 19991 12156
rect 19935 12020 19991 12076
rect 19935 11940 19991 11996
rect 22825 12180 22881 12236
rect 22825 12100 22881 12156
rect 22825 12020 22881 12076
rect 22825 11940 22881 11996
rect 25715 12180 25771 12236
rect 25715 12100 25771 12156
rect 25715 12020 25771 12076
rect 25715 11940 25771 11996
rect 28605 12180 28661 12236
rect 28605 12100 28661 12156
rect 28605 12020 28661 12076
rect 28605 11940 28661 11996
rect 31495 12180 31551 12236
rect 31495 12100 31551 12156
rect 31495 12020 31551 12076
rect 31495 11940 31551 11996
rect 34385 12180 34441 12236
rect 34385 12100 34441 12156
rect 34385 12020 34441 12076
rect 34385 11940 34441 11996
rect 37275 12180 37331 12236
rect 37275 12100 37331 12156
rect 37275 12020 37331 12076
rect 37275 11940 37331 11996
rect 40165 12180 40221 12236
rect 40165 12100 40221 12156
rect 40165 12020 40221 12076
rect 40165 11940 40221 11996
rect 43055 12180 43111 12236
rect 43055 12100 43111 12156
rect 43055 12020 43111 12076
rect 43055 11940 43111 11996
rect 45945 12180 46001 12236
rect 45945 12100 46001 12156
rect 45945 12020 46001 12076
rect 45945 11940 46001 11996
rect 48892 12180 48948 12236
rect 48892 12100 48948 12156
rect 48892 12020 48948 12076
rect 48892 11940 48948 11996
rect 49754 12180 49810 12236
rect 49834 12180 49890 12236
rect 49754 12100 49810 12156
rect 49834 12100 49890 12156
rect 49754 12020 49810 12076
rect 49834 12020 49890 12076
rect 49754 11940 49810 11996
rect 49834 11940 49890 11996
rect 53048 12180 53104 12236
rect 53048 12100 53104 12156
rect 53048 12020 53104 12076
rect 53048 11940 53104 11996
rect 53206 12180 53262 12236
rect 53206 12100 53262 12156
rect 53206 12020 53262 12076
rect 53206 11940 53262 11996
rect 53562 12180 53618 12236
rect 53562 12100 53618 12156
rect 53562 12020 53618 12076
rect 53562 11940 53618 11996
rect 54880 12180 54936 12236
rect 54880 12100 54936 12156
rect 54880 12020 54936 12076
rect 54880 11940 54936 11996
rect 55473 12180 55529 12236
rect 55473 12100 55529 12156
rect 55473 12020 55529 12076
rect 55473 11940 55529 11996
rect 56619 12180 56675 12236
rect 56619 12100 56675 12156
rect 56619 12020 56675 12076
rect 56619 11940 56675 11996
rect 58055 12180 58111 12236
rect 58135 12180 58191 12236
rect 58055 12100 58111 12156
rect 58135 12100 58191 12156
rect 58055 12020 58111 12076
rect 58135 12020 58191 12076
rect 58055 11940 58111 11996
rect 58135 11940 58191 11996
rect 59298 12180 59354 12236
rect 59298 12100 59354 12156
rect 59298 12020 59354 12076
rect 59298 11940 59354 11996
rect 59456 12180 59512 12236
rect 59456 12100 59512 12156
rect 59456 12020 59512 12076
rect 59456 11940 59512 11996
rect 59764 12180 59820 12236
rect 59764 12100 59820 12156
rect 59764 12020 59820 12076
rect 59764 11940 59820 11996
rect 59910 12180 59966 12236
rect 59910 12100 59966 12156
rect 59910 12020 59966 12076
rect 59910 11940 59966 11996
rect 60046 12180 60102 12236
rect 60126 12180 60182 12236
rect 60046 12100 60102 12156
rect 60126 12100 60182 12156
rect 60046 12020 60102 12076
rect 60126 12020 60182 12076
rect 60046 11940 60102 11996
rect 60126 11940 60182 11996
rect 62418 12180 62474 12236
rect 62498 12180 62554 12236
rect 62418 12100 62474 12156
rect 62498 12100 62554 12156
rect 62418 12020 62474 12076
rect 62498 12020 62554 12076
rect 62418 11940 62474 11996
rect 62498 11940 62554 11996
rect 63682 18128 63738 18184
rect 63590 15816 63646 15872
rect 63590 11500 63592 11520
rect 63592 11500 63644 11520
rect 63644 11500 63646 11520
rect 63590 11464 63646 11500
rect 63590 10512 63646 10568
rect 63498 10004 63500 10024
rect 63500 10004 63552 10024
rect 63552 10004 63554 10024
rect 63498 9968 63554 10004
rect 63498 9832 63554 9888
rect 1864 2180 1920 2236
rect 1944 2180 2000 2236
rect 2024 2180 2080 2236
rect 2104 2180 2160 2236
rect 1864 2100 1920 2156
rect 1944 2100 2000 2156
rect 2024 2100 2080 2156
rect 2104 2100 2160 2156
rect 1864 2020 1920 2076
rect 1944 2020 2000 2076
rect 2024 2020 2080 2076
rect 2104 2020 2160 2076
rect 1864 1940 1920 1996
rect 1944 1940 2000 1996
rect 2024 1940 2080 1996
rect 2104 1940 2160 1996
rect 4216 4532 4272 4588
rect 4296 4532 4352 4588
rect 4376 4532 4432 4588
rect 4456 4532 4512 4588
rect 4216 4452 4272 4508
rect 4296 4452 4352 4508
rect 4376 4452 4432 4508
rect 4456 4452 4512 4508
rect 4216 4378 4272 4428
rect 4296 4378 4352 4428
rect 4376 4378 4432 4428
rect 4456 4378 4512 4428
rect 4216 4372 4262 4378
rect 4262 4372 4272 4378
rect 4296 4372 4326 4378
rect 4326 4372 4338 4378
rect 4338 4372 4352 4378
rect 4376 4372 4390 4378
rect 4390 4372 4402 4378
rect 4402 4372 4432 4378
rect 4456 4372 4466 4378
rect 4466 4372 4512 4378
rect 4216 4326 4262 4348
rect 4262 4326 4272 4348
rect 4296 4326 4326 4348
rect 4326 4326 4338 4348
rect 4338 4326 4352 4348
rect 4376 4326 4390 4348
rect 4390 4326 4402 4348
rect 4402 4326 4432 4348
rect 4456 4326 4466 4348
rect 4466 4326 4512 4348
rect 4216 4292 4272 4326
rect 4296 4292 4352 4326
rect 4376 4292 4432 4326
rect 4456 4292 4512 4326
rect 11864 2180 11920 2236
rect 11944 2180 12000 2236
rect 12024 2180 12080 2236
rect 12104 2180 12160 2236
rect 11864 2100 11920 2156
rect 11944 2100 12000 2156
rect 12024 2100 12080 2156
rect 12104 2100 12160 2156
rect 11864 2020 11920 2076
rect 11944 2020 12000 2076
rect 12024 2020 12080 2076
rect 12104 2020 12160 2076
rect 11864 1940 11920 1996
rect 11944 1940 12000 1996
rect 12024 1940 12080 1996
rect 12104 1940 12160 1996
rect 14216 4532 14272 4588
rect 14296 4532 14352 4588
rect 14376 4532 14432 4588
rect 14456 4532 14512 4588
rect 14216 4452 14272 4508
rect 14296 4452 14352 4508
rect 14376 4452 14432 4508
rect 14456 4452 14512 4508
rect 14216 4378 14272 4428
rect 14296 4378 14352 4428
rect 14376 4378 14432 4428
rect 14456 4378 14512 4428
rect 14216 4372 14262 4378
rect 14262 4372 14272 4378
rect 14296 4372 14326 4378
rect 14326 4372 14338 4378
rect 14338 4372 14352 4378
rect 14376 4372 14390 4378
rect 14390 4372 14402 4378
rect 14402 4372 14432 4378
rect 14456 4372 14466 4378
rect 14466 4372 14512 4378
rect 14216 4326 14262 4348
rect 14262 4326 14272 4348
rect 14296 4326 14326 4348
rect 14326 4326 14338 4348
rect 14338 4326 14352 4348
rect 14376 4326 14390 4348
rect 14390 4326 14402 4348
rect 14402 4326 14432 4348
rect 14456 4326 14466 4348
rect 14466 4326 14512 4348
rect 14216 4292 14272 4326
rect 14296 4292 14352 4326
rect 14376 4292 14432 4326
rect 14456 4292 14512 4326
rect 21864 2180 21920 2236
rect 21944 2180 22000 2236
rect 22024 2180 22080 2236
rect 22104 2180 22160 2236
rect 21864 2100 21920 2156
rect 21944 2100 22000 2156
rect 22024 2100 22080 2156
rect 22104 2100 22160 2156
rect 21864 2020 21920 2076
rect 21944 2020 22000 2076
rect 22024 2020 22080 2076
rect 22104 2020 22160 2076
rect 21864 1940 21920 1996
rect 21944 1940 22000 1996
rect 22024 1940 22080 1996
rect 22104 1940 22160 1996
rect 24216 4532 24272 4588
rect 24296 4532 24352 4588
rect 24376 4532 24432 4588
rect 24456 4532 24512 4588
rect 24216 4452 24272 4508
rect 24296 4452 24352 4508
rect 24376 4452 24432 4508
rect 24456 4452 24512 4508
rect 24216 4378 24272 4428
rect 24296 4378 24352 4428
rect 24376 4378 24432 4428
rect 24456 4378 24512 4428
rect 24216 4372 24262 4378
rect 24262 4372 24272 4378
rect 24296 4372 24326 4378
rect 24326 4372 24338 4378
rect 24338 4372 24352 4378
rect 24376 4372 24390 4378
rect 24390 4372 24402 4378
rect 24402 4372 24432 4378
rect 24456 4372 24466 4378
rect 24466 4372 24512 4378
rect 24216 4326 24262 4348
rect 24262 4326 24272 4348
rect 24296 4326 24326 4348
rect 24326 4326 24338 4348
rect 24338 4326 24352 4348
rect 24376 4326 24390 4348
rect 24390 4326 24402 4348
rect 24402 4326 24432 4348
rect 24456 4326 24466 4348
rect 24466 4326 24512 4348
rect 24216 4292 24272 4326
rect 24296 4292 24352 4326
rect 24376 4292 24432 4326
rect 24456 4292 24512 4326
rect 26882 3440 26938 3496
rect 29826 4020 29828 4040
rect 29828 4020 29880 4040
rect 29880 4020 29882 4040
rect 29826 3984 29882 4020
rect 30746 5344 30802 5400
rect 31574 6160 31630 6216
rect 30930 5072 30986 5128
rect 29734 2760 29790 2816
rect 30562 2352 30618 2408
rect 31666 5228 31722 5264
rect 31666 5208 31668 5228
rect 31668 5208 31720 5228
rect 31720 5208 31722 5228
rect 32218 5208 32274 5264
rect 32494 5228 32550 5264
rect 32494 5208 32496 5228
rect 32496 5208 32548 5228
rect 32548 5208 32550 5228
rect 32402 5108 32404 5128
rect 32404 5108 32456 5128
rect 32456 5108 32458 5128
rect 32402 5072 32458 5108
rect 32402 4936 32458 4992
rect 32310 4120 32366 4176
rect 31666 3168 31722 3224
rect 32402 3304 32458 3360
rect 32218 3032 32274 3088
rect 32586 3576 32642 3632
rect 31864 2180 31920 2236
rect 31944 2180 32000 2236
rect 32024 2180 32080 2236
rect 32104 2180 32160 2236
rect 31864 2100 31920 2156
rect 31944 2100 32000 2156
rect 32024 2100 32080 2156
rect 32104 2100 32160 2156
rect 31864 2020 31920 2076
rect 31944 2020 32000 2076
rect 32024 2020 32080 2076
rect 32104 2020 32160 2076
rect 31864 1940 31920 1996
rect 31944 1940 32000 1996
rect 32024 1940 32080 1996
rect 32104 1940 32160 1996
rect 33598 4120 33654 4176
rect 33414 3848 33470 3904
rect 33414 2896 33470 2952
rect 33782 6296 33838 6352
rect 34058 5072 34114 5128
rect 33966 4800 34022 4856
rect 34702 4800 34758 4856
rect 34216 4532 34272 4588
rect 34296 4532 34352 4588
rect 34376 4532 34432 4588
rect 34456 4532 34512 4588
rect 34886 5344 34942 5400
rect 33782 3304 33838 3360
rect 34216 4452 34272 4508
rect 34296 4452 34352 4508
rect 34376 4452 34432 4508
rect 34456 4452 34512 4508
rect 34216 4378 34272 4428
rect 34296 4378 34352 4428
rect 34376 4378 34432 4428
rect 34456 4378 34512 4428
rect 34216 4372 34262 4378
rect 34262 4372 34272 4378
rect 34296 4372 34326 4378
rect 34326 4372 34338 4378
rect 34338 4372 34352 4378
rect 34376 4372 34390 4378
rect 34390 4372 34402 4378
rect 34402 4372 34432 4378
rect 34456 4372 34466 4378
rect 34466 4372 34512 4378
rect 34216 4326 34262 4348
rect 34262 4326 34272 4348
rect 34296 4326 34326 4348
rect 34326 4326 34338 4348
rect 34338 4326 34352 4348
rect 34376 4326 34390 4348
rect 34390 4326 34402 4348
rect 34402 4326 34432 4348
rect 34456 4326 34466 4348
rect 34466 4326 34512 4348
rect 34216 4292 34272 4326
rect 34296 4292 34352 4326
rect 34376 4292 34432 4326
rect 34456 4292 34512 4326
rect 34058 4120 34114 4176
rect 33966 3712 34022 3768
rect 33966 3340 33968 3360
rect 33968 3340 34020 3360
rect 34020 3340 34022 3360
rect 33966 3304 34022 3340
rect 35806 5344 35862 5400
rect 35622 5072 35678 5128
rect 34978 4800 35034 4856
rect 33874 2488 33930 2544
rect 33966 1300 33968 1320
rect 33968 1300 34020 1320
rect 34020 1300 34022 1320
rect 33966 1264 34022 1300
rect 35162 4120 35218 4176
rect 35438 4156 35440 4176
rect 35440 4156 35492 4176
rect 35492 4156 35494 4176
rect 35438 4120 35494 4156
rect 34978 3340 34980 3360
rect 34980 3340 35032 3360
rect 35032 3340 35034 3360
rect 34978 3304 35034 3340
rect 34886 2352 34942 2408
rect 35254 3712 35310 3768
rect 35714 3712 35770 3768
rect 35438 2896 35494 2952
rect 36266 4936 36322 4992
rect 40222 6432 40278 6488
rect 37922 5208 37978 5264
rect 36082 3168 36138 3224
rect 36266 3848 36322 3904
rect 36174 2760 36230 2816
rect 36634 3712 36690 3768
rect 36450 3032 36506 3088
rect 37462 3032 37518 3088
rect 42706 5616 42762 5672
rect 44730 5788 44732 5808
rect 44732 5788 44784 5808
rect 44784 5788 44786 5808
rect 44730 5752 44786 5788
rect 44216 4532 44272 4588
rect 44296 4532 44352 4588
rect 44376 4532 44432 4588
rect 44456 4532 44512 4588
rect 44216 4452 44272 4508
rect 44296 4452 44352 4508
rect 44376 4452 44432 4508
rect 44456 4452 44512 4508
rect 44216 4378 44272 4428
rect 44296 4378 44352 4428
rect 44376 4378 44432 4428
rect 44456 4378 44512 4428
rect 44216 4372 44262 4378
rect 44262 4372 44272 4378
rect 44296 4372 44326 4378
rect 44326 4372 44338 4378
rect 44338 4372 44352 4378
rect 44376 4372 44390 4378
rect 44390 4372 44402 4378
rect 44402 4372 44432 4378
rect 44456 4372 44466 4378
rect 44466 4372 44512 4378
rect 44216 4326 44262 4348
rect 44262 4326 44272 4348
rect 44296 4326 44326 4348
rect 44326 4326 44338 4348
rect 44338 4326 44352 4348
rect 44376 4326 44390 4348
rect 44390 4326 44402 4348
rect 44402 4326 44432 4348
rect 44456 4326 44466 4348
rect 44466 4326 44512 4348
rect 44216 4292 44272 4326
rect 44296 4292 44352 4326
rect 44376 4292 44432 4326
rect 44456 4292 44512 4326
rect 41864 2180 41920 2236
rect 41944 2180 42000 2236
rect 42024 2180 42080 2236
rect 42104 2180 42160 2236
rect 41864 2100 41920 2156
rect 41944 2100 42000 2156
rect 42024 2100 42080 2156
rect 42104 2100 42160 2156
rect 41142 1672 41198 1728
rect 41864 2020 41920 2076
rect 41944 2020 42000 2076
rect 42024 2020 42080 2076
rect 42104 2020 42160 2076
rect 41864 1940 41920 1996
rect 41944 1940 42000 1996
rect 42024 1940 42080 1996
rect 42104 1940 42160 1996
rect 45282 4936 45338 4992
rect 59274 7792 59330 7848
rect 59634 7656 59690 7712
rect 61290 7656 61346 7712
rect 61474 7656 61530 7712
rect 58254 7520 58310 7576
rect 57334 7112 57390 7168
rect 55034 6704 55090 6760
rect 52366 6568 52422 6624
rect 48502 4936 48558 4992
rect 47950 1672 48006 1728
rect 50342 3712 50398 3768
rect 50894 3188 50950 3224
rect 50894 3168 50896 3188
rect 50896 3168 50948 3188
rect 50948 3168 50950 3188
rect 51170 3168 51226 3224
rect 51864 2180 51920 2236
rect 51944 2180 52000 2236
rect 52024 2180 52080 2236
rect 52104 2180 52160 2236
rect 51864 2100 51920 2156
rect 51944 2100 52000 2156
rect 52024 2100 52080 2156
rect 52104 2100 52160 2156
rect 51864 2020 51920 2076
rect 51944 2020 52000 2076
rect 52024 2020 52080 2076
rect 52104 2020 52160 2076
rect 51864 1940 51920 1996
rect 51944 1940 52000 1996
rect 52024 1940 52080 1996
rect 52104 1940 52160 1996
rect 53746 5480 53802 5536
rect 54216 4532 54272 4588
rect 54296 4532 54352 4588
rect 54376 4532 54432 4588
rect 54456 4532 54512 4588
rect 54216 4452 54272 4508
rect 54296 4452 54352 4508
rect 54376 4452 54432 4508
rect 54456 4452 54512 4508
rect 54216 4378 54272 4428
rect 54296 4378 54352 4428
rect 54376 4378 54432 4428
rect 54456 4378 54512 4428
rect 54216 4372 54262 4378
rect 54262 4372 54272 4378
rect 54296 4372 54326 4378
rect 54326 4372 54338 4378
rect 54338 4372 54352 4378
rect 54376 4372 54390 4378
rect 54390 4372 54402 4378
rect 54402 4372 54432 4378
rect 54456 4372 54466 4378
rect 54466 4372 54512 4378
rect 54216 4326 54262 4348
rect 54262 4326 54272 4348
rect 54296 4326 54326 4348
rect 54326 4326 54338 4348
rect 54338 4326 54352 4348
rect 54376 4326 54390 4348
rect 54390 4326 54402 4348
rect 54402 4326 54432 4348
rect 54456 4326 54466 4348
rect 54466 4326 54512 4348
rect 54216 4292 54272 4326
rect 54296 4292 54352 4326
rect 54376 4292 54432 4326
rect 54456 4292 54512 4326
rect 53010 3340 53012 3360
rect 53012 3340 53064 3360
rect 53064 3340 53066 3360
rect 53010 3304 53066 3340
rect 53378 3304 53434 3360
rect 56506 5888 56562 5944
rect 58714 3168 58770 3224
rect 61290 7384 61346 7440
rect 60278 5108 60280 5128
rect 60280 5108 60332 5128
rect 60332 5108 60334 5128
rect 60278 5072 60334 5108
rect 61750 5244 61752 5264
rect 61752 5244 61804 5264
rect 61804 5244 61806 5264
rect 61750 5208 61806 5244
rect 60462 4936 60518 4992
rect 61106 4936 61162 4992
rect 62394 5244 62396 5264
rect 62396 5244 62448 5264
rect 62448 5244 62450 5264
rect 61198 4120 61254 4176
rect 62394 5208 62450 5244
rect 62394 3168 62450 3224
rect 62670 7248 62726 7304
rect 62578 6976 62634 7032
rect 62854 6024 62910 6080
rect 61864 2180 61920 2236
rect 61944 2180 62000 2236
rect 62024 2180 62080 2236
rect 62104 2180 62160 2236
rect 61864 2100 61920 2156
rect 61944 2100 62000 2156
rect 62024 2100 62080 2156
rect 62104 2100 62160 2156
rect 61864 2020 61920 2076
rect 61944 2020 62000 2076
rect 62024 2020 62080 2076
rect 62104 2020 62160 2076
rect 61864 1940 61920 1996
rect 61944 1940 62000 1996
rect 62024 1940 62080 1996
rect 62104 1940 62160 1996
rect 63590 6024 63646 6080
rect 63866 41248 63922 41304
rect 64326 6432 64382 6488
rect 64602 11736 64658 11792
rect 64602 7656 64658 7712
rect 64216 4532 64272 4588
rect 64296 4532 64352 4588
rect 64376 4532 64432 4588
rect 64456 4532 64512 4588
rect 64216 4452 64272 4508
rect 64296 4452 64352 4508
rect 64376 4452 64432 4508
rect 64456 4452 64512 4508
rect 64216 4378 64272 4428
rect 64296 4378 64352 4428
rect 64376 4378 64432 4428
rect 64456 4378 64512 4428
rect 64216 4372 64262 4378
rect 64262 4372 64272 4378
rect 64296 4372 64326 4378
rect 64326 4372 64338 4378
rect 64338 4372 64352 4378
rect 64376 4372 64390 4378
rect 64390 4372 64402 4378
rect 64402 4372 64432 4378
rect 64456 4372 64466 4378
rect 64466 4372 64512 4378
rect 64216 4326 64262 4348
rect 64262 4326 64272 4348
rect 64296 4326 64326 4348
rect 64326 4326 64338 4348
rect 64338 4326 64352 4348
rect 64376 4326 64390 4348
rect 64390 4326 64402 4348
rect 64402 4326 64432 4348
rect 64456 4326 64466 4348
rect 64466 4326 64512 4348
rect 64216 4292 64272 4326
rect 64296 4292 64352 4326
rect 64376 4292 64432 4326
rect 64456 4292 64512 4326
rect 63682 4120 63738 4176
rect 65706 46996 65708 47016
rect 65708 46996 65760 47016
rect 65760 46996 65762 47016
rect 65706 46960 65762 46996
rect 65982 46996 65984 47016
rect 65984 46996 66036 47016
rect 66036 46996 66038 47016
rect 65982 46960 66038 46996
rect 65706 38548 65762 38584
rect 65706 38528 65708 38548
rect 65708 38528 65760 38548
rect 65760 38528 65762 38548
rect 65430 34720 65486 34776
rect 65338 11736 65394 11792
rect 65246 5072 65302 5128
rect 66074 12688 66130 12744
rect 66074 9152 66130 9208
rect 66258 22344 66314 22400
rect 66166 8880 66222 8936
rect 65798 3984 65854 4040
rect 66258 7792 66314 7848
rect 66534 22616 66590 22672
rect 66074 3440 66130 3496
rect 66442 7384 66498 7440
rect 67178 23604 67180 23624
rect 67180 23604 67232 23624
rect 67232 23604 67234 23624
rect 67178 23568 67234 23604
rect 67270 23432 67326 23488
rect 67638 6160 67694 6216
rect 67822 6296 67878 6352
rect 68558 5616 68614 5672
rect 68650 4800 68706 4856
rect 71864 82180 71920 82236
rect 71944 82180 72000 82236
rect 72024 82180 72080 82236
rect 72104 82180 72160 82236
rect 71864 82118 71910 82156
rect 71910 82118 71920 82156
rect 71944 82118 71974 82156
rect 71974 82118 71986 82156
rect 71986 82118 72000 82156
rect 72024 82118 72038 82156
rect 72038 82118 72050 82156
rect 72050 82118 72080 82156
rect 72104 82118 72114 82156
rect 72114 82118 72160 82156
rect 71864 82100 71920 82118
rect 71944 82100 72000 82118
rect 72024 82100 72080 82118
rect 72104 82100 72160 82118
rect 71864 82020 71920 82076
rect 71944 82020 72000 82076
rect 72024 82020 72080 82076
rect 72104 82020 72160 82076
rect 71864 81940 71920 81996
rect 71944 81940 72000 81996
rect 72024 81940 72080 81996
rect 72104 81940 72160 81996
rect 71864 72180 71920 72236
rect 71944 72180 72000 72236
rect 72024 72180 72080 72236
rect 72104 72180 72160 72236
rect 71864 72100 71920 72156
rect 71944 72100 72000 72156
rect 72024 72100 72080 72156
rect 72104 72100 72160 72156
rect 71864 72020 71920 72076
rect 71944 72020 72000 72076
rect 72024 72020 72080 72076
rect 72104 72020 72160 72076
rect 71864 71940 71920 71996
rect 71944 71940 72000 71996
rect 72024 71940 72080 71996
rect 72104 71940 72160 71996
rect 71864 62180 71920 62236
rect 71944 62180 72000 62236
rect 72024 62180 72080 62236
rect 72104 62180 72160 62236
rect 71864 62100 71920 62156
rect 71944 62100 72000 62156
rect 72024 62100 72080 62156
rect 72104 62100 72160 62156
rect 71864 62020 71920 62076
rect 71944 62020 72000 62076
rect 72024 62020 72080 62076
rect 72104 62020 72160 62076
rect 71864 61940 71920 61996
rect 71944 61940 72000 61996
rect 72024 61940 72080 61996
rect 72104 61940 72160 61996
rect 71864 52180 71920 52236
rect 71944 52180 72000 52236
rect 72024 52180 72080 52236
rect 72104 52180 72160 52236
rect 71864 52100 71920 52156
rect 71944 52100 72000 52156
rect 72024 52100 72080 52156
rect 72104 52100 72160 52156
rect 71864 52020 71920 52076
rect 71944 52020 72000 52076
rect 72024 52020 72080 52076
rect 72104 52020 72160 52076
rect 71864 51940 71920 51996
rect 71944 51940 72000 51996
rect 72024 51940 72080 51996
rect 72104 51940 72160 51996
rect 69478 5752 69534 5808
rect 71864 42180 71920 42236
rect 71944 42180 72000 42236
rect 72024 42180 72080 42236
rect 72104 42180 72160 42236
rect 71864 42100 71920 42156
rect 71944 42100 72000 42156
rect 72024 42100 72080 42156
rect 72104 42100 72160 42156
rect 71864 42020 71920 42076
rect 71944 42020 72000 42076
rect 72024 42020 72080 42076
rect 72104 42020 72160 42076
rect 71864 41940 71920 41996
rect 71944 41940 72000 41996
rect 72024 41940 72080 41996
rect 72104 41940 72160 41996
rect 69938 3576 69994 3632
rect 71864 32180 71920 32236
rect 71944 32180 72000 32236
rect 72024 32180 72080 32236
rect 72104 32180 72160 32236
rect 71864 32122 71920 32156
rect 71944 32122 72000 32156
rect 72024 32122 72080 32156
rect 72104 32122 72160 32156
rect 71864 32100 71910 32122
rect 71910 32100 71920 32122
rect 71944 32100 71974 32122
rect 71974 32100 71986 32122
rect 71986 32100 72000 32122
rect 72024 32100 72038 32122
rect 72038 32100 72050 32122
rect 72050 32100 72080 32122
rect 72104 32100 72114 32122
rect 72114 32100 72160 32122
rect 71864 32070 71910 32076
rect 71910 32070 71920 32076
rect 71944 32070 71974 32076
rect 71974 32070 71986 32076
rect 71986 32070 72000 32076
rect 72024 32070 72038 32076
rect 72038 32070 72050 32076
rect 72050 32070 72080 32076
rect 72104 32070 72114 32076
rect 72114 32070 72160 32076
rect 71864 32020 71920 32070
rect 71944 32020 72000 32070
rect 72024 32020 72080 32070
rect 72104 32020 72160 32070
rect 71864 31940 71920 31996
rect 71944 31940 72000 31996
rect 72024 31940 72080 31996
rect 72104 31940 72160 31996
rect 71864 22180 71920 22236
rect 71944 22180 72000 22236
rect 72024 22180 72080 22236
rect 72104 22180 72160 22236
rect 71864 22100 71920 22156
rect 71944 22100 72000 22156
rect 72024 22100 72080 22156
rect 72104 22100 72160 22156
rect 71864 22020 71920 22076
rect 71944 22020 72000 22076
rect 72024 22020 72080 22076
rect 72104 22020 72160 22076
rect 71864 21940 71920 21996
rect 71944 21940 72000 21996
rect 72024 21940 72080 21996
rect 72104 21940 72160 21996
rect 71864 12180 71920 12236
rect 71944 12180 72000 12236
rect 72024 12180 72080 12236
rect 72104 12180 72160 12236
rect 71864 12100 71920 12156
rect 71944 12100 72000 12156
rect 72024 12100 72080 12156
rect 72104 12100 72160 12156
rect 71864 12020 71920 12076
rect 71944 12020 72000 12076
rect 72024 12020 72080 12076
rect 72104 12020 72160 12076
rect 71864 11940 71920 11996
rect 71944 11940 72000 11996
rect 72024 11940 72080 11996
rect 72104 11940 72160 11996
rect 74216 84532 74272 84588
rect 74296 84532 74352 84588
rect 74376 84532 74432 84588
rect 74456 84532 74512 84588
rect 74216 84452 74272 84508
rect 74296 84452 74352 84508
rect 74376 84452 74432 84508
rect 74456 84452 74512 84508
rect 74216 84372 74272 84428
rect 74296 84372 74352 84428
rect 74376 84372 74432 84428
rect 74456 84372 74512 84428
rect 74216 84292 74272 84348
rect 74296 84292 74352 84348
rect 74376 84292 74432 84348
rect 74456 84292 74512 84348
rect 74216 74532 74272 74588
rect 74296 74532 74352 74588
rect 74376 74532 74432 74588
rect 74456 74532 74512 74588
rect 74216 74452 74272 74508
rect 74296 74452 74352 74508
rect 74376 74452 74432 74508
rect 74456 74452 74512 74508
rect 74216 74372 74272 74428
rect 74296 74372 74352 74428
rect 74376 74372 74432 74428
rect 74456 74372 74512 74428
rect 74216 74292 74272 74348
rect 74296 74292 74352 74348
rect 74376 74292 74432 74348
rect 74456 74292 74512 74348
rect 74216 64532 74272 64588
rect 74296 64532 74352 64588
rect 74376 64532 74432 64588
rect 74456 64532 74512 64588
rect 74216 64452 74272 64508
rect 74296 64452 74352 64508
rect 74376 64452 74432 64508
rect 74456 64452 74512 64508
rect 74216 64372 74272 64428
rect 74296 64372 74352 64428
rect 74376 64372 74432 64428
rect 74456 64372 74512 64428
rect 74216 64292 74272 64348
rect 74296 64292 74352 64348
rect 74376 64292 74432 64348
rect 74456 64292 74512 64348
rect 74216 54532 74272 54588
rect 74296 54532 74352 54588
rect 74376 54532 74432 54588
rect 74456 54532 74512 54588
rect 74216 54452 74272 54508
rect 74296 54452 74352 54508
rect 74376 54452 74432 54508
rect 74456 54452 74512 54508
rect 74216 54426 74272 54428
rect 74296 54426 74352 54428
rect 74376 54426 74432 54428
rect 74456 54426 74512 54428
rect 74216 54374 74262 54426
rect 74262 54374 74272 54426
rect 74296 54374 74326 54426
rect 74326 54374 74338 54426
rect 74338 54374 74352 54426
rect 74376 54374 74390 54426
rect 74390 54374 74402 54426
rect 74402 54374 74432 54426
rect 74456 54374 74466 54426
rect 74466 54374 74512 54426
rect 74216 54372 74272 54374
rect 74296 54372 74352 54374
rect 74376 54372 74432 54374
rect 74456 54372 74512 54374
rect 74216 54292 74272 54348
rect 74296 54292 74352 54348
rect 74376 54292 74432 54348
rect 74456 54292 74512 54348
rect 74216 44582 74262 44588
rect 74262 44582 74272 44588
rect 74296 44582 74326 44588
rect 74326 44582 74338 44588
rect 74338 44582 74352 44588
rect 74376 44582 74390 44588
rect 74390 44582 74402 44588
rect 74402 44582 74432 44588
rect 74456 44582 74466 44588
rect 74466 44582 74512 44588
rect 74216 44532 74272 44582
rect 74296 44532 74352 44582
rect 74376 44532 74432 44582
rect 74456 44532 74512 44582
rect 74216 44452 74272 44508
rect 74296 44452 74352 44508
rect 74376 44452 74432 44508
rect 74456 44452 74512 44508
rect 74216 44372 74272 44428
rect 74296 44372 74352 44428
rect 74376 44372 74432 44428
rect 74456 44372 74512 44428
rect 74216 44292 74272 44348
rect 74296 44292 74352 44348
rect 74376 44292 74432 44348
rect 74456 44292 74512 44348
rect 74216 34532 74272 34588
rect 74296 34532 74352 34588
rect 74376 34532 74432 34588
rect 74456 34532 74512 34588
rect 74216 34452 74272 34508
rect 74296 34452 74352 34508
rect 74376 34452 74432 34508
rect 74456 34452 74512 34508
rect 74216 34372 74272 34428
rect 74296 34372 74352 34428
rect 74376 34372 74432 34428
rect 74456 34372 74512 34428
rect 74216 34292 74272 34348
rect 74296 34292 74352 34348
rect 74376 34292 74432 34348
rect 74456 34292 74512 34348
rect 74216 24532 74272 24588
rect 74296 24532 74352 24588
rect 74376 24532 74432 24588
rect 74456 24532 74512 24588
rect 74216 24452 74272 24508
rect 74296 24452 74352 24508
rect 74376 24452 74432 24508
rect 74456 24452 74512 24508
rect 74216 24372 74272 24428
rect 74296 24372 74352 24428
rect 74376 24372 74432 24428
rect 74456 24372 74512 24428
rect 74216 24292 74272 24348
rect 74296 24292 74352 24348
rect 74376 24292 74432 24348
rect 74456 24292 74512 24348
rect 74216 14532 74272 14588
rect 74296 14532 74352 14588
rect 74376 14532 74432 14588
rect 74456 14532 74512 14588
rect 74216 14452 74272 14508
rect 74296 14452 74352 14508
rect 74376 14452 74432 14508
rect 74456 14452 74512 14508
rect 74216 14372 74272 14428
rect 74296 14372 74352 14428
rect 74376 14372 74432 14428
rect 74456 14372 74512 14428
rect 74216 14292 74272 14348
rect 74296 14292 74352 14348
rect 74376 14292 74432 14348
rect 74456 14292 74512 14348
rect 74216 4532 74272 4588
rect 74296 4532 74352 4588
rect 74376 4532 74432 4588
rect 74456 4532 74512 4588
rect 74216 4452 74272 4508
rect 74296 4452 74352 4508
rect 74376 4452 74432 4508
rect 74456 4452 74512 4508
rect 74216 4378 74272 4428
rect 74296 4378 74352 4428
rect 74376 4378 74432 4428
rect 74456 4378 74512 4428
rect 74216 4372 74262 4378
rect 74262 4372 74272 4378
rect 74296 4372 74326 4378
rect 74326 4372 74338 4378
rect 74338 4372 74352 4378
rect 74376 4372 74390 4378
rect 74390 4372 74402 4378
rect 74402 4372 74432 4378
rect 74456 4372 74466 4378
rect 74466 4372 74512 4378
rect 74216 4326 74262 4348
rect 74262 4326 74272 4348
rect 74296 4326 74326 4348
rect 74326 4326 74338 4348
rect 74338 4326 74352 4348
rect 74376 4326 74390 4348
rect 74390 4326 74402 4348
rect 74402 4326 74432 4348
rect 74456 4326 74466 4348
rect 74466 4326 74512 4348
rect 74216 4292 74272 4326
rect 74296 4292 74352 4326
rect 74376 4292 74432 4326
rect 74456 4292 74512 4326
rect 71864 2180 71920 2236
rect 71944 2180 72000 2236
rect 72024 2180 72080 2236
rect 72104 2180 72160 2236
rect 71864 2100 71920 2156
rect 71944 2100 72000 2156
rect 72024 2100 72080 2156
rect 72104 2100 72160 2156
rect 71864 2020 71920 2076
rect 71944 2020 72000 2076
rect 72024 2020 72080 2076
rect 72104 2020 72160 2076
rect 71864 1940 71920 1996
rect 71944 1940 72000 1996
rect 72024 1940 72080 1996
rect 72104 1940 72160 1996
<< metal3 >>
rect 964 84592 75028 84616
rect 964 84588 4740 84592
rect 964 84532 2136 84588
rect 2192 84532 4740 84588
rect 964 84528 4740 84532
rect 4804 84528 4820 84592
rect 4884 84528 4900 84592
rect 4964 84528 4980 84592
rect 5044 84528 5060 84592
rect 5124 84528 5140 84592
rect 5204 84528 5220 84592
rect 5284 84588 10740 84592
rect 5284 84532 5632 84588
rect 5688 84532 8522 84588
rect 8578 84532 10740 84588
rect 5284 84528 10740 84532
rect 10804 84528 10820 84592
rect 10884 84528 10900 84592
rect 10964 84528 10980 84592
rect 11044 84528 11060 84592
rect 11124 84528 11140 84592
rect 11204 84528 11220 84592
rect 11284 84588 16740 84592
rect 11284 84532 11412 84588
rect 11468 84532 14302 84588
rect 14358 84532 16740 84588
rect 11284 84528 16740 84532
rect 16804 84528 16820 84592
rect 16884 84528 16900 84592
rect 16964 84528 16980 84592
rect 17044 84528 17060 84592
rect 17124 84528 17140 84592
rect 17204 84588 17220 84592
rect 17284 84588 22740 84592
rect 17284 84532 20082 84588
rect 20138 84532 22740 84588
rect 17204 84528 17220 84532
rect 17284 84528 22740 84532
rect 22804 84528 22820 84592
rect 22884 84528 22900 84592
rect 22964 84588 22980 84592
rect 22964 84532 22972 84588
rect 22964 84528 22980 84532
rect 23044 84528 23060 84592
rect 23124 84528 23140 84592
rect 23204 84528 23220 84592
rect 23284 84588 28740 84592
rect 28804 84588 28820 84592
rect 23284 84532 25862 84588
rect 25918 84532 28740 84588
rect 28808 84532 28820 84588
rect 23284 84528 28740 84532
rect 28804 84528 28820 84532
rect 28884 84528 28900 84592
rect 28964 84528 28980 84592
rect 29044 84528 29060 84592
rect 29124 84528 29140 84592
rect 29204 84528 29220 84592
rect 29284 84588 34740 84592
rect 29284 84532 31642 84588
rect 31698 84532 34532 84588
rect 34588 84532 34740 84588
rect 29284 84528 34740 84532
rect 34804 84528 34820 84592
rect 34884 84528 34900 84592
rect 34964 84528 34980 84592
rect 35044 84528 35060 84592
rect 35124 84528 35140 84592
rect 35204 84528 35220 84592
rect 35284 84588 40740 84592
rect 35284 84532 37422 84588
rect 37478 84532 40312 84588
rect 40368 84532 40740 84588
rect 35284 84528 40740 84532
rect 40804 84528 40820 84592
rect 40884 84528 40900 84592
rect 40964 84528 40980 84592
rect 41044 84528 41060 84592
rect 41124 84528 41140 84592
rect 41204 84528 41220 84592
rect 41284 84588 46740 84592
rect 41284 84532 43202 84588
rect 43258 84532 46092 84588
rect 46148 84532 46740 84588
rect 41284 84528 46740 84532
rect 46804 84528 46820 84592
rect 46884 84528 46900 84592
rect 46964 84528 46980 84592
rect 47044 84528 47060 84592
rect 47124 84528 47140 84592
rect 47204 84528 47220 84592
rect 47284 84588 52740 84592
rect 47284 84532 49100 84588
rect 49156 84532 52329 84588
rect 52385 84532 52740 84588
rect 47284 84528 52740 84532
rect 52804 84528 52820 84592
rect 52884 84528 52900 84592
rect 52964 84528 52980 84592
rect 53044 84528 53060 84592
rect 53124 84528 53140 84592
rect 53204 84528 53220 84592
rect 53284 84588 58740 84592
rect 53284 84532 53730 84588
rect 53786 84532 53898 84588
rect 53954 84532 54642 84588
rect 54698 84532 55032 84588
rect 55088 84532 55748 84588
rect 55804 84532 56326 84588
rect 56382 84532 56771 84588
rect 56827 84532 57075 84588
rect 57131 84532 57917 84588
rect 57973 84532 58557 84588
rect 58613 84532 58740 84588
rect 53284 84528 58740 84532
rect 58804 84528 58820 84592
rect 58884 84528 58900 84592
rect 58964 84528 58980 84592
rect 59044 84528 59060 84592
rect 59124 84528 59140 84592
rect 59204 84528 59220 84592
rect 59284 84588 64740 84592
rect 59284 84532 60418 84588
rect 60474 84532 60576 84588
rect 60632 84532 62620 84588
rect 62676 84532 62700 84588
rect 62756 84532 64740 84588
rect 59284 84528 64740 84532
rect 64804 84528 64820 84592
rect 64884 84528 64900 84592
rect 64964 84528 64980 84592
rect 65044 84528 65060 84592
rect 65124 84528 65140 84592
rect 65204 84528 65220 84592
rect 65284 84528 70740 84592
rect 70804 84528 70820 84592
rect 70884 84528 70900 84592
rect 70964 84528 70980 84592
rect 71044 84528 71060 84592
rect 71124 84528 71140 84592
rect 71204 84528 71220 84592
rect 71284 84588 75028 84592
rect 71284 84532 74216 84588
rect 74272 84532 74296 84588
rect 74352 84532 74376 84588
rect 74432 84532 74456 84588
rect 74512 84532 75028 84588
rect 71284 84528 75028 84532
rect 964 84512 75028 84528
rect 964 84508 4740 84512
rect 964 84452 2136 84508
rect 2192 84452 4740 84508
rect 964 84448 4740 84452
rect 4804 84448 4820 84512
rect 4884 84448 4900 84512
rect 4964 84448 4980 84512
rect 5044 84448 5060 84512
rect 5124 84448 5140 84512
rect 5204 84448 5220 84512
rect 5284 84508 10740 84512
rect 5284 84452 5632 84508
rect 5688 84452 8522 84508
rect 8578 84452 10740 84508
rect 5284 84448 10740 84452
rect 10804 84448 10820 84512
rect 10884 84448 10900 84512
rect 10964 84448 10980 84512
rect 11044 84448 11060 84512
rect 11124 84448 11140 84512
rect 11204 84448 11220 84512
rect 11284 84508 16740 84512
rect 11284 84452 11412 84508
rect 11468 84452 14302 84508
rect 14358 84452 16740 84508
rect 11284 84448 16740 84452
rect 16804 84448 16820 84512
rect 16884 84448 16900 84512
rect 16964 84448 16980 84512
rect 17044 84448 17060 84512
rect 17124 84448 17140 84512
rect 17204 84508 17220 84512
rect 17284 84508 22740 84512
rect 17284 84452 20082 84508
rect 20138 84452 22740 84508
rect 17204 84448 17220 84452
rect 17284 84448 22740 84452
rect 22804 84448 22820 84512
rect 22884 84448 22900 84512
rect 22964 84508 22980 84512
rect 22964 84452 22972 84508
rect 22964 84448 22980 84452
rect 23044 84448 23060 84512
rect 23124 84448 23140 84512
rect 23204 84448 23220 84512
rect 23284 84508 28740 84512
rect 28804 84508 28820 84512
rect 23284 84452 25862 84508
rect 25918 84452 28740 84508
rect 28808 84452 28820 84508
rect 23284 84448 28740 84452
rect 28804 84448 28820 84452
rect 28884 84448 28900 84512
rect 28964 84448 28980 84512
rect 29044 84448 29060 84512
rect 29124 84448 29140 84512
rect 29204 84448 29220 84512
rect 29284 84508 34740 84512
rect 29284 84452 31642 84508
rect 31698 84452 34532 84508
rect 34588 84452 34740 84508
rect 29284 84448 34740 84452
rect 34804 84448 34820 84512
rect 34884 84448 34900 84512
rect 34964 84448 34980 84512
rect 35044 84448 35060 84512
rect 35124 84448 35140 84512
rect 35204 84448 35220 84512
rect 35284 84508 40740 84512
rect 35284 84452 37422 84508
rect 37478 84452 40312 84508
rect 40368 84452 40740 84508
rect 35284 84448 40740 84452
rect 40804 84448 40820 84512
rect 40884 84448 40900 84512
rect 40964 84448 40980 84512
rect 41044 84448 41060 84512
rect 41124 84448 41140 84512
rect 41204 84448 41220 84512
rect 41284 84508 46740 84512
rect 41284 84452 43202 84508
rect 43258 84452 46092 84508
rect 46148 84452 46740 84508
rect 41284 84448 46740 84452
rect 46804 84448 46820 84512
rect 46884 84448 46900 84512
rect 46964 84448 46980 84512
rect 47044 84448 47060 84512
rect 47124 84448 47140 84512
rect 47204 84448 47220 84512
rect 47284 84508 52740 84512
rect 47284 84452 49100 84508
rect 49156 84452 52329 84508
rect 52385 84452 52740 84508
rect 47284 84448 52740 84452
rect 52804 84448 52820 84512
rect 52884 84448 52900 84512
rect 52964 84448 52980 84512
rect 53044 84448 53060 84512
rect 53124 84448 53140 84512
rect 53204 84448 53220 84512
rect 53284 84508 58740 84512
rect 53284 84452 53730 84508
rect 53786 84452 53898 84508
rect 53954 84452 54642 84508
rect 54698 84452 55032 84508
rect 55088 84452 55748 84508
rect 55804 84452 56326 84508
rect 56382 84452 56771 84508
rect 56827 84452 57075 84508
rect 57131 84452 57917 84508
rect 57973 84452 58557 84508
rect 58613 84452 58740 84508
rect 53284 84448 58740 84452
rect 58804 84448 58820 84512
rect 58884 84448 58900 84512
rect 58964 84448 58980 84512
rect 59044 84448 59060 84512
rect 59124 84448 59140 84512
rect 59204 84448 59220 84512
rect 59284 84508 64740 84512
rect 59284 84452 60418 84508
rect 60474 84452 60576 84508
rect 60632 84452 62620 84508
rect 62676 84452 62700 84508
rect 62756 84452 64740 84508
rect 59284 84448 64740 84452
rect 64804 84448 64820 84512
rect 64884 84448 64900 84512
rect 64964 84448 64980 84512
rect 65044 84448 65060 84512
rect 65124 84448 65140 84512
rect 65204 84448 65220 84512
rect 65284 84448 70740 84512
rect 70804 84448 70820 84512
rect 70884 84448 70900 84512
rect 70964 84448 70980 84512
rect 71044 84448 71060 84512
rect 71124 84448 71140 84512
rect 71204 84448 71220 84512
rect 71284 84508 75028 84512
rect 71284 84452 74216 84508
rect 74272 84452 74296 84508
rect 74352 84452 74376 84508
rect 74432 84452 74456 84508
rect 74512 84452 75028 84508
rect 71284 84448 75028 84452
rect 964 84432 75028 84448
rect 964 84428 4740 84432
rect 964 84372 2136 84428
rect 2192 84372 4740 84428
rect 964 84368 4740 84372
rect 4804 84368 4820 84432
rect 4884 84368 4900 84432
rect 4964 84368 4980 84432
rect 5044 84368 5060 84432
rect 5124 84368 5140 84432
rect 5204 84368 5220 84432
rect 5284 84428 10740 84432
rect 5284 84372 5632 84428
rect 5688 84372 8522 84428
rect 8578 84372 10740 84428
rect 5284 84368 10740 84372
rect 10804 84368 10820 84432
rect 10884 84368 10900 84432
rect 10964 84368 10980 84432
rect 11044 84368 11060 84432
rect 11124 84368 11140 84432
rect 11204 84368 11220 84432
rect 11284 84428 16740 84432
rect 11284 84372 11412 84428
rect 11468 84372 14302 84428
rect 14358 84372 16740 84428
rect 11284 84368 16740 84372
rect 16804 84368 16820 84432
rect 16884 84368 16900 84432
rect 16964 84368 16980 84432
rect 17044 84368 17060 84432
rect 17124 84368 17140 84432
rect 17204 84428 17220 84432
rect 17284 84428 22740 84432
rect 17284 84372 20082 84428
rect 20138 84372 22740 84428
rect 17204 84368 17220 84372
rect 17284 84368 22740 84372
rect 22804 84368 22820 84432
rect 22884 84368 22900 84432
rect 22964 84428 22980 84432
rect 22964 84372 22972 84428
rect 22964 84368 22980 84372
rect 23044 84368 23060 84432
rect 23124 84368 23140 84432
rect 23204 84368 23220 84432
rect 23284 84428 28740 84432
rect 28804 84428 28820 84432
rect 23284 84372 25862 84428
rect 25918 84372 28740 84428
rect 28808 84372 28820 84428
rect 23284 84368 28740 84372
rect 28804 84368 28820 84372
rect 28884 84368 28900 84432
rect 28964 84368 28980 84432
rect 29044 84368 29060 84432
rect 29124 84368 29140 84432
rect 29204 84368 29220 84432
rect 29284 84428 34740 84432
rect 29284 84372 31642 84428
rect 31698 84372 34532 84428
rect 34588 84372 34740 84428
rect 29284 84368 34740 84372
rect 34804 84368 34820 84432
rect 34884 84368 34900 84432
rect 34964 84368 34980 84432
rect 35044 84368 35060 84432
rect 35124 84368 35140 84432
rect 35204 84368 35220 84432
rect 35284 84428 40740 84432
rect 35284 84372 37422 84428
rect 37478 84372 40312 84428
rect 40368 84372 40740 84428
rect 35284 84368 40740 84372
rect 40804 84368 40820 84432
rect 40884 84368 40900 84432
rect 40964 84368 40980 84432
rect 41044 84368 41060 84432
rect 41124 84368 41140 84432
rect 41204 84368 41220 84432
rect 41284 84428 46740 84432
rect 41284 84372 43202 84428
rect 43258 84372 46092 84428
rect 46148 84372 46740 84428
rect 41284 84368 46740 84372
rect 46804 84368 46820 84432
rect 46884 84368 46900 84432
rect 46964 84368 46980 84432
rect 47044 84368 47060 84432
rect 47124 84368 47140 84432
rect 47204 84368 47220 84432
rect 47284 84428 52740 84432
rect 47284 84372 49100 84428
rect 49156 84372 52329 84428
rect 52385 84372 52740 84428
rect 47284 84368 52740 84372
rect 52804 84368 52820 84432
rect 52884 84368 52900 84432
rect 52964 84368 52980 84432
rect 53044 84368 53060 84432
rect 53124 84368 53140 84432
rect 53204 84368 53220 84432
rect 53284 84428 58740 84432
rect 53284 84372 53730 84428
rect 53786 84372 53898 84428
rect 53954 84372 54642 84428
rect 54698 84372 55032 84428
rect 55088 84372 55748 84428
rect 55804 84372 56326 84428
rect 56382 84372 56771 84428
rect 56827 84372 57075 84428
rect 57131 84372 57917 84428
rect 57973 84372 58557 84428
rect 58613 84372 58740 84428
rect 53284 84368 58740 84372
rect 58804 84368 58820 84432
rect 58884 84368 58900 84432
rect 58964 84368 58980 84432
rect 59044 84368 59060 84432
rect 59124 84368 59140 84432
rect 59204 84368 59220 84432
rect 59284 84428 64740 84432
rect 59284 84372 60418 84428
rect 60474 84372 60576 84428
rect 60632 84372 62620 84428
rect 62676 84372 62700 84428
rect 62756 84372 64740 84428
rect 59284 84368 64740 84372
rect 64804 84368 64820 84432
rect 64884 84368 64900 84432
rect 64964 84368 64980 84432
rect 65044 84368 65060 84432
rect 65124 84368 65140 84432
rect 65204 84368 65220 84432
rect 65284 84368 70740 84432
rect 70804 84368 70820 84432
rect 70884 84368 70900 84432
rect 70964 84368 70980 84432
rect 71044 84368 71060 84432
rect 71124 84368 71140 84432
rect 71204 84368 71220 84432
rect 71284 84428 75028 84432
rect 71284 84372 74216 84428
rect 74272 84372 74296 84428
rect 74352 84372 74376 84428
rect 74432 84372 74456 84428
rect 74512 84372 75028 84428
rect 71284 84368 75028 84372
rect 964 84352 75028 84368
rect 964 84348 4740 84352
rect 964 84292 2136 84348
rect 2192 84292 4740 84348
rect 964 84288 4740 84292
rect 4804 84288 4820 84352
rect 4884 84288 4900 84352
rect 4964 84288 4980 84352
rect 5044 84288 5060 84352
rect 5124 84288 5140 84352
rect 5204 84288 5220 84352
rect 5284 84348 10740 84352
rect 5284 84292 5632 84348
rect 5688 84292 8522 84348
rect 8578 84292 10740 84348
rect 5284 84288 10740 84292
rect 10804 84288 10820 84352
rect 10884 84288 10900 84352
rect 10964 84288 10980 84352
rect 11044 84288 11060 84352
rect 11124 84288 11140 84352
rect 11204 84288 11220 84352
rect 11284 84348 16740 84352
rect 11284 84292 11412 84348
rect 11468 84292 14302 84348
rect 14358 84292 16740 84348
rect 11284 84288 16740 84292
rect 16804 84288 16820 84352
rect 16884 84288 16900 84352
rect 16964 84288 16980 84352
rect 17044 84288 17060 84352
rect 17124 84288 17140 84352
rect 17204 84348 17220 84352
rect 17284 84348 22740 84352
rect 17284 84292 20082 84348
rect 20138 84292 22740 84348
rect 17204 84288 17220 84292
rect 17284 84288 22740 84292
rect 22804 84288 22820 84352
rect 22884 84288 22900 84352
rect 22964 84348 22980 84352
rect 22964 84292 22972 84348
rect 22964 84288 22980 84292
rect 23044 84288 23060 84352
rect 23124 84288 23140 84352
rect 23204 84288 23220 84352
rect 23284 84348 28740 84352
rect 28804 84348 28820 84352
rect 23284 84292 25862 84348
rect 25918 84292 28740 84348
rect 28808 84292 28820 84348
rect 23284 84288 28740 84292
rect 28804 84288 28820 84292
rect 28884 84288 28900 84352
rect 28964 84288 28980 84352
rect 29044 84288 29060 84352
rect 29124 84288 29140 84352
rect 29204 84288 29220 84352
rect 29284 84348 34740 84352
rect 29284 84292 31642 84348
rect 31698 84292 34532 84348
rect 34588 84292 34740 84348
rect 29284 84288 34740 84292
rect 34804 84288 34820 84352
rect 34884 84288 34900 84352
rect 34964 84288 34980 84352
rect 35044 84288 35060 84352
rect 35124 84288 35140 84352
rect 35204 84288 35220 84352
rect 35284 84348 40740 84352
rect 35284 84292 37422 84348
rect 37478 84292 40312 84348
rect 40368 84292 40740 84348
rect 35284 84288 40740 84292
rect 40804 84288 40820 84352
rect 40884 84288 40900 84352
rect 40964 84288 40980 84352
rect 41044 84288 41060 84352
rect 41124 84288 41140 84352
rect 41204 84288 41220 84352
rect 41284 84348 46740 84352
rect 41284 84292 43202 84348
rect 43258 84292 46092 84348
rect 46148 84292 46740 84348
rect 41284 84288 46740 84292
rect 46804 84288 46820 84352
rect 46884 84288 46900 84352
rect 46964 84288 46980 84352
rect 47044 84288 47060 84352
rect 47124 84288 47140 84352
rect 47204 84288 47220 84352
rect 47284 84348 52740 84352
rect 47284 84292 49100 84348
rect 49156 84292 52329 84348
rect 52385 84292 52740 84348
rect 47284 84288 52740 84292
rect 52804 84288 52820 84352
rect 52884 84288 52900 84352
rect 52964 84288 52980 84352
rect 53044 84288 53060 84352
rect 53124 84288 53140 84352
rect 53204 84288 53220 84352
rect 53284 84348 58740 84352
rect 53284 84292 53730 84348
rect 53786 84292 53898 84348
rect 53954 84292 54642 84348
rect 54698 84292 55032 84348
rect 55088 84292 55748 84348
rect 55804 84292 56326 84348
rect 56382 84292 56771 84348
rect 56827 84292 57075 84348
rect 57131 84292 57917 84348
rect 57973 84292 58557 84348
rect 58613 84292 58740 84348
rect 53284 84288 58740 84292
rect 58804 84288 58820 84352
rect 58884 84288 58900 84352
rect 58964 84288 58980 84352
rect 59044 84288 59060 84352
rect 59124 84288 59140 84352
rect 59204 84288 59220 84352
rect 59284 84348 64740 84352
rect 59284 84292 60418 84348
rect 60474 84292 60576 84348
rect 60632 84292 62620 84348
rect 62676 84292 62700 84348
rect 62756 84292 64740 84348
rect 59284 84288 64740 84292
rect 64804 84288 64820 84352
rect 64884 84288 64900 84352
rect 64964 84288 64980 84352
rect 65044 84288 65060 84352
rect 65124 84288 65140 84352
rect 65204 84288 65220 84352
rect 65284 84288 70740 84352
rect 70804 84288 70820 84352
rect 70884 84288 70900 84352
rect 70964 84288 70980 84352
rect 71044 84288 71060 84352
rect 71124 84288 71140 84352
rect 71204 84288 71220 84352
rect 71284 84348 75028 84352
rect 71284 84292 74216 84348
rect 74272 84292 74296 84348
rect 74352 84292 74376 84348
rect 74432 84292 74456 84348
rect 74512 84292 75028 84348
rect 71284 84288 75028 84292
rect 964 84264 75028 84288
rect 964 82240 75028 82264
rect 964 82176 1740 82240
rect 1804 82176 1820 82240
rect 1884 82176 1900 82240
rect 1964 82176 1980 82240
rect 2044 82176 2060 82240
rect 2124 82176 2140 82240
rect 2204 82176 2220 82240
rect 2284 82236 7740 82240
rect 2332 82180 2356 82236
rect 2412 82180 5485 82236
rect 5541 82180 7740 82236
rect 2284 82176 7740 82180
rect 7804 82176 7820 82240
rect 7884 82176 7900 82240
rect 7964 82176 7980 82240
rect 8044 82176 8060 82240
rect 8124 82176 8140 82240
rect 8204 82176 8220 82240
rect 8284 82236 13740 82240
rect 8284 82180 8375 82236
rect 8431 82180 11265 82236
rect 11321 82180 13740 82236
rect 8284 82176 13740 82180
rect 13804 82176 13820 82240
rect 13884 82176 13900 82240
rect 13964 82176 13980 82240
rect 14044 82176 14060 82240
rect 14124 82176 14140 82240
rect 14204 82236 14220 82240
rect 14211 82180 14220 82236
rect 14204 82176 14220 82180
rect 14284 82236 19740 82240
rect 14284 82180 17045 82236
rect 17101 82180 19740 82236
rect 14284 82176 19740 82180
rect 19804 82176 19820 82240
rect 19884 82176 19900 82240
rect 19964 82236 19980 82240
rect 19964 82176 19980 82180
rect 20044 82176 20060 82240
rect 20124 82176 20140 82240
rect 20204 82176 20220 82240
rect 20284 82236 25740 82240
rect 20284 82180 22825 82236
rect 22881 82180 25715 82236
rect 20284 82176 25740 82180
rect 25804 82176 25820 82240
rect 25884 82176 25900 82240
rect 25964 82176 25980 82240
rect 26044 82176 26060 82240
rect 26124 82176 26140 82240
rect 26204 82176 26220 82240
rect 26284 82236 31740 82240
rect 26284 82180 28605 82236
rect 28661 82180 31495 82236
rect 31551 82180 31740 82236
rect 26284 82176 31740 82180
rect 31804 82176 31820 82240
rect 31884 82176 31900 82240
rect 31964 82176 31980 82240
rect 32044 82176 32060 82240
rect 32124 82176 32140 82240
rect 32204 82176 32220 82240
rect 32284 82236 37740 82240
rect 32284 82180 34385 82236
rect 34441 82180 37275 82236
rect 37331 82180 37740 82236
rect 32284 82176 37740 82180
rect 37804 82176 37820 82240
rect 37884 82176 37900 82240
rect 37964 82176 37980 82240
rect 38044 82176 38060 82240
rect 38124 82176 38140 82240
rect 38204 82176 38220 82240
rect 38284 82236 43740 82240
rect 38284 82180 40165 82236
rect 40221 82180 43055 82236
rect 43111 82180 43740 82236
rect 38284 82176 43740 82180
rect 43804 82176 43820 82240
rect 43884 82176 43900 82240
rect 43964 82176 43980 82240
rect 44044 82176 44060 82240
rect 44124 82176 44140 82240
rect 44204 82176 44220 82240
rect 44284 82236 49740 82240
rect 49804 82236 49820 82240
rect 49884 82236 49900 82240
rect 44284 82180 45945 82236
rect 46001 82180 48892 82236
rect 48948 82180 49740 82236
rect 49810 82180 49820 82236
rect 49890 82180 49900 82236
rect 44284 82176 49740 82180
rect 49804 82176 49820 82180
rect 49884 82176 49900 82180
rect 49964 82176 49980 82240
rect 50044 82176 50060 82240
rect 50124 82176 50140 82240
rect 50204 82176 50220 82240
rect 50284 82236 55740 82240
rect 50284 82180 53048 82236
rect 53104 82180 53206 82236
rect 53262 82180 53562 82236
rect 53618 82180 54880 82236
rect 54936 82180 55473 82236
rect 55529 82180 55740 82236
rect 50284 82176 55740 82180
rect 55804 82176 55820 82240
rect 55884 82176 55900 82240
rect 55964 82176 55980 82240
rect 56044 82176 56060 82240
rect 56124 82176 56140 82240
rect 56204 82176 56220 82240
rect 56284 82236 61740 82240
rect 56284 82180 56619 82236
rect 56675 82180 58055 82236
rect 58111 82180 58135 82236
rect 58191 82180 59298 82236
rect 59354 82180 59456 82236
rect 59512 82180 59764 82236
rect 59820 82180 59910 82236
rect 59966 82180 60046 82236
rect 60102 82180 60126 82236
rect 60182 82180 61740 82236
rect 56284 82176 61740 82180
rect 61804 82176 61820 82240
rect 61884 82176 61900 82240
rect 61964 82176 61980 82240
rect 62044 82176 62060 82240
rect 62124 82176 62140 82240
rect 62204 82176 62220 82240
rect 62284 82236 67740 82240
rect 62284 82180 62418 82236
rect 62474 82180 62498 82236
rect 62554 82180 67740 82236
rect 62284 82176 67740 82180
rect 67804 82176 67820 82240
rect 67884 82176 67900 82240
rect 67964 82176 67980 82240
rect 68044 82176 68060 82240
rect 68124 82176 68140 82240
rect 68204 82176 68220 82240
rect 68284 82236 73740 82240
rect 68284 82180 71864 82236
rect 71920 82180 71944 82236
rect 72000 82180 72024 82236
rect 72080 82180 72104 82236
rect 72160 82180 73740 82236
rect 68284 82176 73740 82180
rect 73804 82176 73820 82240
rect 73884 82176 73900 82240
rect 73964 82176 73980 82240
rect 74044 82176 74060 82240
rect 74124 82176 74140 82240
rect 74204 82176 74220 82240
rect 74284 82176 75028 82240
rect 964 82160 75028 82176
rect 964 82096 1740 82160
rect 1804 82096 1820 82160
rect 1884 82096 1900 82160
rect 1964 82096 1980 82160
rect 2044 82096 2060 82160
rect 2124 82096 2140 82160
rect 2204 82096 2220 82160
rect 2284 82156 7740 82160
rect 2332 82100 2356 82156
rect 2412 82100 5485 82156
rect 5541 82100 7740 82156
rect 2284 82096 7740 82100
rect 7804 82096 7820 82160
rect 7884 82096 7900 82160
rect 7964 82096 7980 82160
rect 8044 82096 8060 82160
rect 8124 82096 8140 82160
rect 8204 82096 8220 82160
rect 8284 82156 13740 82160
rect 8284 82100 8375 82156
rect 8431 82100 11265 82156
rect 11321 82100 13740 82156
rect 8284 82096 13740 82100
rect 13804 82096 13820 82160
rect 13884 82096 13900 82160
rect 13964 82096 13980 82160
rect 14044 82096 14060 82160
rect 14124 82096 14140 82160
rect 14204 82156 14220 82160
rect 14211 82100 14220 82156
rect 14204 82096 14220 82100
rect 14284 82156 19740 82160
rect 14284 82100 17045 82156
rect 17101 82100 19740 82156
rect 14284 82096 19740 82100
rect 19804 82096 19820 82160
rect 19884 82096 19900 82160
rect 19964 82156 19980 82160
rect 19964 82096 19980 82100
rect 20044 82096 20060 82160
rect 20124 82096 20140 82160
rect 20204 82096 20220 82160
rect 20284 82156 25740 82160
rect 20284 82100 22825 82156
rect 22881 82100 25715 82156
rect 20284 82096 25740 82100
rect 25804 82096 25820 82160
rect 25884 82096 25900 82160
rect 25964 82096 25980 82160
rect 26044 82096 26060 82160
rect 26124 82096 26140 82160
rect 26204 82096 26220 82160
rect 26284 82156 31740 82160
rect 26284 82100 28605 82156
rect 28661 82100 31495 82156
rect 31551 82100 31740 82156
rect 26284 82096 31740 82100
rect 31804 82096 31820 82160
rect 31884 82096 31900 82160
rect 31964 82096 31980 82160
rect 32044 82096 32060 82160
rect 32124 82096 32140 82160
rect 32204 82096 32220 82160
rect 32284 82156 37740 82160
rect 32284 82100 34385 82156
rect 34441 82100 37275 82156
rect 37331 82100 37740 82156
rect 32284 82096 37740 82100
rect 37804 82096 37820 82160
rect 37884 82096 37900 82160
rect 37964 82096 37980 82160
rect 38044 82096 38060 82160
rect 38124 82096 38140 82160
rect 38204 82096 38220 82160
rect 38284 82156 43740 82160
rect 38284 82100 40165 82156
rect 40221 82100 43055 82156
rect 43111 82100 43740 82156
rect 38284 82096 43740 82100
rect 43804 82096 43820 82160
rect 43884 82096 43900 82160
rect 43964 82096 43980 82160
rect 44044 82096 44060 82160
rect 44124 82096 44140 82160
rect 44204 82096 44220 82160
rect 44284 82156 49740 82160
rect 49804 82156 49820 82160
rect 49884 82156 49900 82160
rect 44284 82100 45945 82156
rect 46001 82100 48892 82156
rect 48948 82100 49740 82156
rect 49810 82100 49820 82156
rect 49890 82100 49900 82156
rect 44284 82096 49740 82100
rect 49804 82096 49820 82100
rect 49884 82096 49900 82100
rect 49964 82096 49980 82160
rect 50044 82096 50060 82160
rect 50124 82096 50140 82160
rect 50204 82096 50220 82160
rect 50284 82156 55740 82160
rect 50284 82100 53048 82156
rect 53104 82100 53206 82156
rect 53262 82100 53562 82156
rect 53618 82100 54880 82156
rect 54936 82100 55473 82156
rect 55529 82100 55740 82156
rect 50284 82096 55740 82100
rect 55804 82096 55820 82160
rect 55884 82096 55900 82160
rect 55964 82096 55980 82160
rect 56044 82096 56060 82160
rect 56124 82096 56140 82160
rect 56204 82096 56220 82160
rect 56284 82156 61740 82160
rect 56284 82100 56619 82156
rect 56675 82100 58055 82156
rect 58111 82100 58135 82156
rect 58191 82100 59298 82156
rect 59354 82100 59456 82156
rect 59512 82100 59764 82156
rect 59820 82100 59910 82156
rect 59966 82100 60046 82156
rect 60102 82100 60126 82156
rect 60182 82100 61740 82156
rect 56284 82096 61740 82100
rect 61804 82096 61820 82160
rect 61884 82096 61900 82160
rect 61964 82096 61980 82160
rect 62044 82096 62060 82160
rect 62124 82096 62140 82160
rect 62204 82096 62220 82160
rect 62284 82156 67740 82160
rect 62284 82100 62418 82156
rect 62474 82100 62498 82156
rect 62554 82100 67740 82156
rect 62284 82096 67740 82100
rect 67804 82096 67820 82160
rect 67884 82096 67900 82160
rect 67964 82096 67980 82160
rect 68044 82096 68060 82160
rect 68124 82096 68140 82160
rect 68204 82096 68220 82160
rect 68284 82156 73740 82160
rect 68284 82100 71864 82156
rect 71920 82100 71944 82156
rect 72000 82100 72024 82156
rect 72080 82100 72104 82156
rect 72160 82100 73740 82156
rect 68284 82096 73740 82100
rect 73804 82096 73820 82160
rect 73884 82096 73900 82160
rect 73964 82096 73980 82160
rect 74044 82096 74060 82160
rect 74124 82096 74140 82160
rect 74204 82096 74220 82160
rect 74284 82096 75028 82160
rect 964 82080 75028 82096
rect 964 82016 1740 82080
rect 1804 82016 1820 82080
rect 1884 82016 1900 82080
rect 1964 82016 1980 82080
rect 2044 82016 2060 82080
rect 2124 82016 2140 82080
rect 2204 82016 2220 82080
rect 2284 82076 7740 82080
rect 2332 82020 2356 82076
rect 2412 82020 5485 82076
rect 5541 82020 7740 82076
rect 2284 82016 7740 82020
rect 7804 82016 7820 82080
rect 7884 82016 7900 82080
rect 7964 82016 7980 82080
rect 8044 82016 8060 82080
rect 8124 82016 8140 82080
rect 8204 82016 8220 82080
rect 8284 82076 13740 82080
rect 8284 82020 8375 82076
rect 8431 82020 11265 82076
rect 11321 82020 13740 82076
rect 8284 82016 13740 82020
rect 13804 82016 13820 82080
rect 13884 82016 13900 82080
rect 13964 82016 13980 82080
rect 14044 82016 14060 82080
rect 14124 82016 14140 82080
rect 14204 82076 14220 82080
rect 14211 82020 14220 82076
rect 14204 82016 14220 82020
rect 14284 82076 19740 82080
rect 14284 82020 17045 82076
rect 17101 82020 19740 82076
rect 14284 82016 19740 82020
rect 19804 82016 19820 82080
rect 19884 82016 19900 82080
rect 19964 82076 19980 82080
rect 19964 82016 19980 82020
rect 20044 82016 20060 82080
rect 20124 82016 20140 82080
rect 20204 82016 20220 82080
rect 20284 82076 25740 82080
rect 20284 82020 22825 82076
rect 22881 82020 25715 82076
rect 20284 82016 25740 82020
rect 25804 82016 25820 82080
rect 25884 82016 25900 82080
rect 25964 82016 25980 82080
rect 26044 82016 26060 82080
rect 26124 82016 26140 82080
rect 26204 82016 26220 82080
rect 26284 82076 31740 82080
rect 26284 82020 28605 82076
rect 28661 82020 31495 82076
rect 31551 82020 31740 82076
rect 26284 82016 31740 82020
rect 31804 82016 31820 82080
rect 31884 82016 31900 82080
rect 31964 82016 31980 82080
rect 32044 82016 32060 82080
rect 32124 82016 32140 82080
rect 32204 82016 32220 82080
rect 32284 82076 37740 82080
rect 32284 82020 34385 82076
rect 34441 82020 37275 82076
rect 37331 82020 37740 82076
rect 32284 82016 37740 82020
rect 37804 82016 37820 82080
rect 37884 82016 37900 82080
rect 37964 82016 37980 82080
rect 38044 82016 38060 82080
rect 38124 82016 38140 82080
rect 38204 82016 38220 82080
rect 38284 82076 43740 82080
rect 38284 82020 40165 82076
rect 40221 82020 43055 82076
rect 43111 82020 43740 82076
rect 38284 82016 43740 82020
rect 43804 82016 43820 82080
rect 43884 82016 43900 82080
rect 43964 82016 43980 82080
rect 44044 82016 44060 82080
rect 44124 82016 44140 82080
rect 44204 82016 44220 82080
rect 44284 82076 49740 82080
rect 49804 82076 49820 82080
rect 49884 82076 49900 82080
rect 44284 82020 45945 82076
rect 46001 82020 48892 82076
rect 48948 82020 49740 82076
rect 49810 82020 49820 82076
rect 49890 82020 49900 82076
rect 44284 82016 49740 82020
rect 49804 82016 49820 82020
rect 49884 82016 49900 82020
rect 49964 82016 49980 82080
rect 50044 82016 50060 82080
rect 50124 82016 50140 82080
rect 50204 82016 50220 82080
rect 50284 82076 55740 82080
rect 50284 82020 53048 82076
rect 53104 82020 53206 82076
rect 53262 82020 53562 82076
rect 53618 82020 54880 82076
rect 54936 82020 55473 82076
rect 55529 82020 55740 82076
rect 50284 82016 55740 82020
rect 55804 82016 55820 82080
rect 55884 82016 55900 82080
rect 55964 82016 55980 82080
rect 56044 82016 56060 82080
rect 56124 82016 56140 82080
rect 56204 82016 56220 82080
rect 56284 82076 61740 82080
rect 56284 82020 56619 82076
rect 56675 82020 58055 82076
rect 58111 82020 58135 82076
rect 58191 82020 59298 82076
rect 59354 82020 59456 82076
rect 59512 82020 59764 82076
rect 59820 82020 59910 82076
rect 59966 82020 60046 82076
rect 60102 82020 60126 82076
rect 60182 82020 61740 82076
rect 56284 82016 61740 82020
rect 61804 82016 61820 82080
rect 61884 82016 61900 82080
rect 61964 82016 61980 82080
rect 62044 82016 62060 82080
rect 62124 82016 62140 82080
rect 62204 82016 62220 82080
rect 62284 82076 67740 82080
rect 62284 82020 62418 82076
rect 62474 82020 62498 82076
rect 62554 82020 67740 82076
rect 62284 82016 67740 82020
rect 67804 82016 67820 82080
rect 67884 82016 67900 82080
rect 67964 82016 67980 82080
rect 68044 82016 68060 82080
rect 68124 82016 68140 82080
rect 68204 82016 68220 82080
rect 68284 82076 73740 82080
rect 68284 82020 71864 82076
rect 71920 82020 71944 82076
rect 72000 82020 72024 82076
rect 72080 82020 72104 82076
rect 72160 82020 73740 82076
rect 68284 82016 73740 82020
rect 73804 82016 73820 82080
rect 73884 82016 73900 82080
rect 73964 82016 73980 82080
rect 74044 82016 74060 82080
rect 74124 82016 74140 82080
rect 74204 82016 74220 82080
rect 74284 82016 75028 82080
rect 964 82000 75028 82016
rect 964 81936 1740 82000
rect 1804 81936 1820 82000
rect 1884 81936 1900 82000
rect 1964 81936 1980 82000
rect 2044 81936 2060 82000
rect 2124 81936 2140 82000
rect 2204 81936 2220 82000
rect 2284 81996 7740 82000
rect 2332 81940 2356 81996
rect 2412 81940 5485 81996
rect 5541 81940 7740 81996
rect 2284 81936 7740 81940
rect 7804 81936 7820 82000
rect 7884 81936 7900 82000
rect 7964 81936 7980 82000
rect 8044 81936 8060 82000
rect 8124 81936 8140 82000
rect 8204 81936 8220 82000
rect 8284 81996 13740 82000
rect 8284 81940 8375 81996
rect 8431 81940 11265 81996
rect 11321 81940 13740 81996
rect 8284 81936 13740 81940
rect 13804 81936 13820 82000
rect 13884 81936 13900 82000
rect 13964 81936 13980 82000
rect 14044 81936 14060 82000
rect 14124 81936 14140 82000
rect 14204 81996 14220 82000
rect 14211 81940 14220 81996
rect 14204 81936 14220 81940
rect 14284 81996 19740 82000
rect 14284 81940 17045 81996
rect 17101 81940 19740 81996
rect 14284 81936 19740 81940
rect 19804 81936 19820 82000
rect 19884 81936 19900 82000
rect 19964 81996 19980 82000
rect 19964 81936 19980 81940
rect 20044 81936 20060 82000
rect 20124 81936 20140 82000
rect 20204 81936 20220 82000
rect 20284 81996 25740 82000
rect 20284 81940 22825 81996
rect 22881 81940 25715 81996
rect 20284 81936 25740 81940
rect 25804 81936 25820 82000
rect 25884 81936 25900 82000
rect 25964 81936 25980 82000
rect 26044 81936 26060 82000
rect 26124 81936 26140 82000
rect 26204 81936 26220 82000
rect 26284 81996 31740 82000
rect 26284 81940 28605 81996
rect 28661 81940 31495 81996
rect 31551 81940 31740 81996
rect 26284 81936 31740 81940
rect 31804 81936 31820 82000
rect 31884 81936 31900 82000
rect 31964 81936 31980 82000
rect 32044 81936 32060 82000
rect 32124 81936 32140 82000
rect 32204 81936 32220 82000
rect 32284 81996 37740 82000
rect 32284 81940 34385 81996
rect 34441 81940 37275 81996
rect 37331 81940 37740 81996
rect 32284 81936 37740 81940
rect 37804 81936 37820 82000
rect 37884 81936 37900 82000
rect 37964 81936 37980 82000
rect 38044 81936 38060 82000
rect 38124 81936 38140 82000
rect 38204 81936 38220 82000
rect 38284 81996 43740 82000
rect 38284 81940 40165 81996
rect 40221 81940 43055 81996
rect 43111 81940 43740 81996
rect 38284 81936 43740 81940
rect 43804 81936 43820 82000
rect 43884 81936 43900 82000
rect 43964 81936 43980 82000
rect 44044 81936 44060 82000
rect 44124 81936 44140 82000
rect 44204 81936 44220 82000
rect 44284 81996 49740 82000
rect 49804 81996 49820 82000
rect 49884 81996 49900 82000
rect 44284 81940 45945 81996
rect 46001 81940 48892 81996
rect 48948 81940 49740 81996
rect 49810 81940 49820 81996
rect 49890 81940 49900 81996
rect 44284 81936 49740 81940
rect 49804 81936 49820 81940
rect 49884 81936 49900 81940
rect 49964 81936 49980 82000
rect 50044 81936 50060 82000
rect 50124 81936 50140 82000
rect 50204 81936 50220 82000
rect 50284 81996 55740 82000
rect 50284 81940 53048 81996
rect 53104 81940 53206 81996
rect 53262 81940 53562 81996
rect 53618 81940 54880 81996
rect 54936 81940 55473 81996
rect 55529 81940 55740 81996
rect 50284 81936 55740 81940
rect 55804 81936 55820 82000
rect 55884 81936 55900 82000
rect 55964 81936 55980 82000
rect 56044 81936 56060 82000
rect 56124 81936 56140 82000
rect 56204 81936 56220 82000
rect 56284 81996 61740 82000
rect 56284 81940 56619 81996
rect 56675 81940 58055 81996
rect 58111 81940 58135 81996
rect 58191 81940 59298 81996
rect 59354 81940 59456 81996
rect 59512 81940 59764 81996
rect 59820 81940 59910 81996
rect 59966 81940 60046 81996
rect 60102 81940 60126 81996
rect 60182 81940 61740 81996
rect 56284 81936 61740 81940
rect 61804 81936 61820 82000
rect 61884 81936 61900 82000
rect 61964 81936 61980 82000
rect 62044 81936 62060 82000
rect 62124 81936 62140 82000
rect 62204 81936 62220 82000
rect 62284 81996 67740 82000
rect 62284 81940 62418 81996
rect 62474 81940 62498 81996
rect 62554 81940 67740 81996
rect 62284 81936 67740 81940
rect 67804 81936 67820 82000
rect 67884 81936 67900 82000
rect 67964 81936 67980 82000
rect 68044 81936 68060 82000
rect 68124 81936 68140 82000
rect 68204 81936 68220 82000
rect 68284 81996 73740 82000
rect 68284 81940 71864 81996
rect 71920 81940 71944 81996
rect 72000 81940 72024 81996
rect 72080 81940 72104 81996
rect 72160 81940 73740 81996
rect 68284 81936 73740 81940
rect 73804 81936 73820 82000
rect 73884 81936 73900 82000
rect 73964 81936 73980 82000
rect 74044 81936 74060 82000
rect 74124 81936 74140 82000
rect 74204 81936 74220 82000
rect 74284 81936 75028 82000
rect 964 81912 75028 81936
rect 964 74592 75028 74616
rect 964 74588 4740 74592
rect 964 74532 2136 74588
rect 2192 74532 4740 74588
rect 964 74528 4740 74532
rect 4804 74528 4820 74592
rect 4884 74528 4900 74592
rect 4964 74528 4980 74592
rect 5044 74528 5060 74592
rect 5124 74528 5140 74592
rect 5204 74528 5220 74592
rect 5284 74588 10740 74592
rect 5284 74532 5632 74588
rect 5688 74532 8522 74588
rect 8578 74532 10740 74588
rect 5284 74528 10740 74532
rect 10804 74528 10820 74592
rect 10884 74528 10900 74592
rect 10964 74528 10980 74592
rect 11044 74528 11060 74592
rect 11124 74528 11140 74592
rect 11204 74528 11220 74592
rect 11284 74588 16740 74592
rect 11284 74532 11412 74588
rect 11468 74532 14302 74588
rect 14358 74532 16740 74588
rect 11284 74528 16740 74532
rect 16804 74528 16820 74592
rect 16884 74528 16900 74592
rect 16964 74528 16980 74592
rect 17044 74528 17060 74592
rect 17124 74528 17140 74592
rect 17204 74588 17220 74592
rect 17284 74588 22740 74592
rect 17284 74532 20082 74588
rect 20138 74532 22740 74588
rect 17204 74528 17220 74532
rect 17284 74528 22740 74532
rect 22804 74528 22820 74592
rect 22884 74528 22900 74592
rect 22964 74588 22980 74592
rect 22964 74532 22972 74588
rect 22964 74528 22980 74532
rect 23044 74528 23060 74592
rect 23124 74528 23140 74592
rect 23204 74528 23220 74592
rect 23284 74588 28740 74592
rect 28804 74588 28820 74592
rect 23284 74532 25862 74588
rect 25918 74532 28740 74588
rect 28808 74532 28820 74588
rect 23284 74528 28740 74532
rect 28804 74528 28820 74532
rect 28884 74528 28900 74592
rect 28964 74528 28980 74592
rect 29044 74528 29060 74592
rect 29124 74528 29140 74592
rect 29204 74528 29220 74592
rect 29284 74588 34740 74592
rect 29284 74532 31642 74588
rect 31698 74532 34532 74588
rect 34588 74532 34740 74588
rect 29284 74528 34740 74532
rect 34804 74528 34820 74592
rect 34884 74528 34900 74592
rect 34964 74528 34980 74592
rect 35044 74528 35060 74592
rect 35124 74528 35140 74592
rect 35204 74528 35220 74592
rect 35284 74588 40740 74592
rect 35284 74532 37422 74588
rect 37478 74532 40312 74588
rect 40368 74532 40740 74588
rect 35284 74528 40740 74532
rect 40804 74528 40820 74592
rect 40884 74528 40900 74592
rect 40964 74528 40980 74592
rect 41044 74528 41060 74592
rect 41124 74528 41140 74592
rect 41204 74528 41220 74592
rect 41284 74588 46740 74592
rect 41284 74532 43202 74588
rect 43258 74532 46092 74588
rect 46148 74532 46740 74588
rect 41284 74528 46740 74532
rect 46804 74528 46820 74592
rect 46884 74528 46900 74592
rect 46964 74528 46980 74592
rect 47044 74528 47060 74592
rect 47124 74528 47140 74592
rect 47204 74528 47220 74592
rect 47284 74588 52740 74592
rect 47284 74532 49100 74588
rect 49156 74532 52329 74588
rect 52385 74532 52740 74588
rect 47284 74528 52740 74532
rect 52804 74528 52820 74592
rect 52884 74528 52900 74592
rect 52964 74528 52980 74592
rect 53044 74528 53060 74592
rect 53124 74528 53140 74592
rect 53204 74528 53220 74592
rect 53284 74588 58740 74592
rect 53284 74532 53730 74588
rect 53786 74532 53898 74588
rect 53954 74532 54642 74588
rect 54698 74532 55032 74588
rect 55088 74532 55748 74588
rect 55804 74532 56326 74588
rect 56382 74532 56771 74588
rect 56827 74532 57075 74588
rect 57131 74532 57917 74588
rect 57973 74532 58557 74588
rect 58613 74532 58740 74588
rect 53284 74528 58740 74532
rect 58804 74528 58820 74592
rect 58884 74528 58900 74592
rect 58964 74528 58980 74592
rect 59044 74528 59060 74592
rect 59124 74528 59140 74592
rect 59204 74528 59220 74592
rect 59284 74588 64740 74592
rect 59284 74532 60418 74588
rect 60474 74532 60576 74588
rect 60632 74532 62620 74588
rect 62676 74532 62700 74588
rect 62756 74532 64740 74588
rect 59284 74528 64740 74532
rect 64804 74528 64820 74592
rect 64884 74528 64900 74592
rect 64964 74528 64980 74592
rect 65044 74528 65060 74592
rect 65124 74528 65140 74592
rect 65204 74528 65220 74592
rect 65284 74528 70740 74592
rect 70804 74528 70820 74592
rect 70884 74528 70900 74592
rect 70964 74528 70980 74592
rect 71044 74528 71060 74592
rect 71124 74528 71140 74592
rect 71204 74528 71220 74592
rect 71284 74588 75028 74592
rect 71284 74532 74216 74588
rect 74272 74532 74296 74588
rect 74352 74532 74376 74588
rect 74432 74532 74456 74588
rect 74512 74532 75028 74588
rect 71284 74528 75028 74532
rect 964 74512 75028 74528
rect 964 74508 4740 74512
rect 964 74452 2136 74508
rect 2192 74452 4740 74508
rect 964 74448 4740 74452
rect 4804 74448 4820 74512
rect 4884 74448 4900 74512
rect 4964 74448 4980 74512
rect 5044 74448 5060 74512
rect 5124 74448 5140 74512
rect 5204 74448 5220 74512
rect 5284 74508 10740 74512
rect 5284 74452 5632 74508
rect 5688 74452 8522 74508
rect 8578 74452 10740 74508
rect 5284 74448 10740 74452
rect 10804 74448 10820 74512
rect 10884 74448 10900 74512
rect 10964 74448 10980 74512
rect 11044 74448 11060 74512
rect 11124 74448 11140 74512
rect 11204 74448 11220 74512
rect 11284 74508 16740 74512
rect 11284 74452 11412 74508
rect 11468 74452 14302 74508
rect 14358 74452 16740 74508
rect 11284 74448 16740 74452
rect 16804 74448 16820 74512
rect 16884 74448 16900 74512
rect 16964 74448 16980 74512
rect 17044 74448 17060 74512
rect 17124 74448 17140 74512
rect 17204 74508 17220 74512
rect 17284 74508 22740 74512
rect 17284 74452 20082 74508
rect 20138 74452 22740 74508
rect 17204 74448 17220 74452
rect 17284 74448 22740 74452
rect 22804 74448 22820 74512
rect 22884 74448 22900 74512
rect 22964 74508 22980 74512
rect 22964 74452 22972 74508
rect 22964 74448 22980 74452
rect 23044 74448 23060 74512
rect 23124 74448 23140 74512
rect 23204 74448 23220 74512
rect 23284 74508 28740 74512
rect 28804 74508 28820 74512
rect 23284 74452 25862 74508
rect 25918 74452 28740 74508
rect 28808 74452 28820 74508
rect 23284 74448 28740 74452
rect 28804 74448 28820 74452
rect 28884 74448 28900 74512
rect 28964 74448 28980 74512
rect 29044 74448 29060 74512
rect 29124 74448 29140 74512
rect 29204 74448 29220 74512
rect 29284 74508 34740 74512
rect 29284 74452 31642 74508
rect 31698 74452 34532 74508
rect 34588 74452 34740 74508
rect 29284 74448 34740 74452
rect 34804 74448 34820 74512
rect 34884 74448 34900 74512
rect 34964 74448 34980 74512
rect 35044 74448 35060 74512
rect 35124 74448 35140 74512
rect 35204 74448 35220 74512
rect 35284 74508 40740 74512
rect 35284 74452 37422 74508
rect 37478 74452 40312 74508
rect 40368 74452 40740 74508
rect 35284 74448 40740 74452
rect 40804 74448 40820 74512
rect 40884 74448 40900 74512
rect 40964 74448 40980 74512
rect 41044 74448 41060 74512
rect 41124 74448 41140 74512
rect 41204 74448 41220 74512
rect 41284 74508 46740 74512
rect 41284 74452 43202 74508
rect 43258 74452 46092 74508
rect 46148 74452 46740 74508
rect 41284 74448 46740 74452
rect 46804 74448 46820 74512
rect 46884 74448 46900 74512
rect 46964 74448 46980 74512
rect 47044 74448 47060 74512
rect 47124 74448 47140 74512
rect 47204 74448 47220 74512
rect 47284 74508 52740 74512
rect 47284 74452 49100 74508
rect 49156 74452 52329 74508
rect 52385 74452 52740 74508
rect 47284 74448 52740 74452
rect 52804 74448 52820 74512
rect 52884 74448 52900 74512
rect 52964 74448 52980 74512
rect 53044 74448 53060 74512
rect 53124 74448 53140 74512
rect 53204 74448 53220 74512
rect 53284 74508 58740 74512
rect 53284 74452 53730 74508
rect 53786 74452 53898 74508
rect 53954 74452 54642 74508
rect 54698 74452 55032 74508
rect 55088 74452 55748 74508
rect 55804 74452 56326 74508
rect 56382 74452 56771 74508
rect 56827 74452 57075 74508
rect 57131 74452 57917 74508
rect 57973 74452 58557 74508
rect 58613 74452 58740 74508
rect 53284 74448 58740 74452
rect 58804 74448 58820 74512
rect 58884 74448 58900 74512
rect 58964 74448 58980 74512
rect 59044 74448 59060 74512
rect 59124 74448 59140 74512
rect 59204 74448 59220 74512
rect 59284 74508 64740 74512
rect 59284 74452 60418 74508
rect 60474 74452 60576 74508
rect 60632 74452 62620 74508
rect 62676 74452 62700 74508
rect 62756 74452 64740 74508
rect 59284 74448 64740 74452
rect 64804 74448 64820 74512
rect 64884 74448 64900 74512
rect 64964 74448 64980 74512
rect 65044 74448 65060 74512
rect 65124 74448 65140 74512
rect 65204 74448 65220 74512
rect 65284 74448 70740 74512
rect 70804 74448 70820 74512
rect 70884 74448 70900 74512
rect 70964 74448 70980 74512
rect 71044 74448 71060 74512
rect 71124 74448 71140 74512
rect 71204 74448 71220 74512
rect 71284 74508 75028 74512
rect 71284 74452 74216 74508
rect 74272 74452 74296 74508
rect 74352 74452 74376 74508
rect 74432 74452 74456 74508
rect 74512 74452 75028 74508
rect 71284 74448 75028 74452
rect 964 74432 75028 74448
rect 964 74428 4740 74432
rect 964 74372 2136 74428
rect 2192 74372 4740 74428
rect 964 74368 4740 74372
rect 4804 74368 4820 74432
rect 4884 74368 4900 74432
rect 4964 74368 4980 74432
rect 5044 74368 5060 74432
rect 5124 74368 5140 74432
rect 5204 74368 5220 74432
rect 5284 74428 10740 74432
rect 5284 74372 5632 74428
rect 5688 74372 8522 74428
rect 8578 74372 10740 74428
rect 5284 74368 10740 74372
rect 10804 74368 10820 74432
rect 10884 74368 10900 74432
rect 10964 74368 10980 74432
rect 11044 74368 11060 74432
rect 11124 74368 11140 74432
rect 11204 74368 11220 74432
rect 11284 74428 16740 74432
rect 11284 74372 11412 74428
rect 11468 74372 14302 74428
rect 14358 74372 16740 74428
rect 11284 74368 16740 74372
rect 16804 74368 16820 74432
rect 16884 74368 16900 74432
rect 16964 74368 16980 74432
rect 17044 74368 17060 74432
rect 17124 74368 17140 74432
rect 17204 74428 17220 74432
rect 17284 74428 22740 74432
rect 17284 74372 20082 74428
rect 20138 74372 22740 74428
rect 17204 74368 17220 74372
rect 17284 74368 22740 74372
rect 22804 74368 22820 74432
rect 22884 74368 22900 74432
rect 22964 74428 22980 74432
rect 22964 74372 22972 74428
rect 22964 74368 22980 74372
rect 23044 74368 23060 74432
rect 23124 74368 23140 74432
rect 23204 74368 23220 74432
rect 23284 74428 28740 74432
rect 28804 74428 28820 74432
rect 23284 74372 25862 74428
rect 25918 74372 28740 74428
rect 28808 74372 28820 74428
rect 23284 74368 28740 74372
rect 28804 74368 28820 74372
rect 28884 74368 28900 74432
rect 28964 74368 28980 74432
rect 29044 74368 29060 74432
rect 29124 74368 29140 74432
rect 29204 74368 29220 74432
rect 29284 74428 34740 74432
rect 29284 74372 31642 74428
rect 31698 74372 34532 74428
rect 34588 74372 34740 74428
rect 29284 74368 34740 74372
rect 34804 74368 34820 74432
rect 34884 74368 34900 74432
rect 34964 74368 34980 74432
rect 35044 74368 35060 74432
rect 35124 74368 35140 74432
rect 35204 74368 35220 74432
rect 35284 74428 40740 74432
rect 35284 74372 37422 74428
rect 37478 74372 40312 74428
rect 40368 74372 40740 74428
rect 35284 74368 40740 74372
rect 40804 74368 40820 74432
rect 40884 74368 40900 74432
rect 40964 74368 40980 74432
rect 41044 74368 41060 74432
rect 41124 74368 41140 74432
rect 41204 74368 41220 74432
rect 41284 74428 46740 74432
rect 41284 74372 43202 74428
rect 43258 74372 46092 74428
rect 46148 74372 46740 74428
rect 41284 74368 46740 74372
rect 46804 74368 46820 74432
rect 46884 74368 46900 74432
rect 46964 74368 46980 74432
rect 47044 74368 47060 74432
rect 47124 74368 47140 74432
rect 47204 74368 47220 74432
rect 47284 74428 52740 74432
rect 47284 74372 49100 74428
rect 49156 74372 52329 74428
rect 52385 74372 52740 74428
rect 47284 74368 52740 74372
rect 52804 74368 52820 74432
rect 52884 74368 52900 74432
rect 52964 74368 52980 74432
rect 53044 74368 53060 74432
rect 53124 74368 53140 74432
rect 53204 74368 53220 74432
rect 53284 74428 58740 74432
rect 53284 74372 53730 74428
rect 53786 74372 53898 74428
rect 53954 74372 54642 74428
rect 54698 74372 55032 74428
rect 55088 74372 55748 74428
rect 55804 74372 56326 74428
rect 56382 74372 56771 74428
rect 56827 74372 57075 74428
rect 57131 74372 57917 74428
rect 57973 74372 58557 74428
rect 58613 74372 58740 74428
rect 53284 74368 58740 74372
rect 58804 74368 58820 74432
rect 58884 74368 58900 74432
rect 58964 74368 58980 74432
rect 59044 74368 59060 74432
rect 59124 74368 59140 74432
rect 59204 74368 59220 74432
rect 59284 74428 64740 74432
rect 59284 74372 60418 74428
rect 60474 74372 60576 74428
rect 60632 74372 62620 74428
rect 62676 74372 62700 74428
rect 62756 74372 64740 74428
rect 59284 74368 64740 74372
rect 64804 74368 64820 74432
rect 64884 74368 64900 74432
rect 64964 74368 64980 74432
rect 65044 74368 65060 74432
rect 65124 74368 65140 74432
rect 65204 74368 65220 74432
rect 65284 74368 70740 74432
rect 70804 74368 70820 74432
rect 70884 74368 70900 74432
rect 70964 74368 70980 74432
rect 71044 74368 71060 74432
rect 71124 74368 71140 74432
rect 71204 74368 71220 74432
rect 71284 74428 75028 74432
rect 71284 74372 74216 74428
rect 74272 74372 74296 74428
rect 74352 74372 74376 74428
rect 74432 74372 74456 74428
rect 74512 74372 75028 74428
rect 71284 74368 75028 74372
rect 964 74352 75028 74368
rect 964 74348 4740 74352
rect 964 74292 2136 74348
rect 2192 74292 4740 74348
rect 964 74288 4740 74292
rect 4804 74288 4820 74352
rect 4884 74288 4900 74352
rect 4964 74288 4980 74352
rect 5044 74288 5060 74352
rect 5124 74288 5140 74352
rect 5204 74288 5220 74352
rect 5284 74348 10740 74352
rect 5284 74292 5632 74348
rect 5688 74292 8522 74348
rect 8578 74292 10740 74348
rect 5284 74288 10740 74292
rect 10804 74288 10820 74352
rect 10884 74288 10900 74352
rect 10964 74288 10980 74352
rect 11044 74288 11060 74352
rect 11124 74288 11140 74352
rect 11204 74288 11220 74352
rect 11284 74348 16740 74352
rect 11284 74292 11412 74348
rect 11468 74292 14302 74348
rect 14358 74292 16740 74348
rect 11284 74288 16740 74292
rect 16804 74288 16820 74352
rect 16884 74288 16900 74352
rect 16964 74288 16980 74352
rect 17044 74288 17060 74352
rect 17124 74288 17140 74352
rect 17204 74348 17220 74352
rect 17284 74348 22740 74352
rect 17284 74292 20082 74348
rect 20138 74292 22740 74348
rect 17204 74288 17220 74292
rect 17284 74288 22740 74292
rect 22804 74288 22820 74352
rect 22884 74288 22900 74352
rect 22964 74348 22980 74352
rect 22964 74292 22972 74348
rect 22964 74288 22980 74292
rect 23044 74288 23060 74352
rect 23124 74288 23140 74352
rect 23204 74288 23220 74352
rect 23284 74348 28740 74352
rect 28804 74348 28820 74352
rect 23284 74292 25862 74348
rect 25918 74292 28740 74348
rect 28808 74292 28820 74348
rect 23284 74288 28740 74292
rect 28804 74288 28820 74292
rect 28884 74288 28900 74352
rect 28964 74288 28980 74352
rect 29044 74288 29060 74352
rect 29124 74288 29140 74352
rect 29204 74288 29220 74352
rect 29284 74348 34740 74352
rect 29284 74292 31642 74348
rect 31698 74292 34532 74348
rect 34588 74292 34740 74348
rect 29284 74288 34740 74292
rect 34804 74288 34820 74352
rect 34884 74288 34900 74352
rect 34964 74288 34980 74352
rect 35044 74288 35060 74352
rect 35124 74288 35140 74352
rect 35204 74288 35220 74352
rect 35284 74348 40740 74352
rect 35284 74292 37422 74348
rect 37478 74292 40312 74348
rect 40368 74292 40740 74348
rect 35284 74288 40740 74292
rect 40804 74288 40820 74352
rect 40884 74288 40900 74352
rect 40964 74288 40980 74352
rect 41044 74288 41060 74352
rect 41124 74288 41140 74352
rect 41204 74288 41220 74352
rect 41284 74348 46740 74352
rect 41284 74292 43202 74348
rect 43258 74292 46092 74348
rect 46148 74292 46740 74348
rect 41284 74288 46740 74292
rect 46804 74288 46820 74352
rect 46884 74288 46900 74352
rect 46964 74288 46980 74352
rect 47044 74288 47060 74352
rect 47124 74288 47140 74352
rect 47204 74288 47220 74352
rect 47284 74348 52740 74352
rect 47284 74292 49100 74348
rect 49156 74292 52329 74348
rect 52385 74292 52740 74348
rect 47284 74288 52740 74292
rect 52804 74288 52820 74352
rect 52884 74288 52900 74352
rect 52964 74288 52980 74352
rect 53044 74288 53060 74352
rect 53124 74288 53140 74352
rect 53204 74288 53220 74352
rect 53284 74348 58740 74352
rect 53284 74292 53730 74348
rect 53786 74292 53898 74348
rect 53954 74292 54642 74348
rect 54698 74292 55032 74348
rect 55088 74292 55748 74348
rect 55804 74292 56326 74348
rect 56382 74292 56771 74348
rect 56827 74292 57075 74348
rect 57131 74292 57917 74348
rect 57973 74292 58557 74348
rect 58613 74292 58740 74348
rect 53284 74288 58740 74292
rect 58804 74288 58820 74352
rect 58884 74288 58900 74352
rect 58964 74288 58980 74352
rect 59044 74288 59060 74352
rect 59124 74288 59140 74352
rect 59204 74288 59220 74352
rect 59284 74348 64740 74352
rect 59284 74292 60418 74348
rect 60474 74292 60576 74348
rect 60632 74292 62620 74348
rect 62676 74292 62700 74348
rect 62756 74292 64740 74348
rect 59284 74288 64740 74292
rect 64804 74288 64820 74352
rect 64884 74288 64900 74352
rect 64964 74288 64980 74352
rect 65044 74288 65060 74352
rect 65124 74288 65140 74352
rect 65204 74288 65220 74352
rect 65284 74288 70740 74352
rect 70804 74288 70820 74352
rect 70884 74288 70900 74352
rect 70964 74288 70980 74352
rect 71044 74288 71060 74352
rect 71124 74288 71140 74352
rect 71204 74288 71220 74352
rect 71284 74348 75028 74352
rect 71284 74292 74216 74348
rect 74272 74292 74296 74348
rect 74352 74292 74376 74348
rect 74432 74292 74456 74348
rect 74512 74292 75028 74348
rect 71284 74288 75028 74292
rect 964 74264 75028 74288
rect 964 72240 75028 72264
rect 964 72176 1740 72240
rect 1804 72176 1820 72240
rect 1884 72176 1900 72240
rect 1964 72176 1980 72240
rect 2044 72176 2060 72240
rect 2124 72176 2140 72240
rect 2204 72176 2220 72240
rect 2284 72236 7740 72240
rect 2332 72180 2356 72236
rect 2412 72180 5485 72236
rect 5541 72180 7740 72236
rect 2284 72176 7740 72180
rect 7804 72176 7820 72240
rect 7884 72176 7900 72240
rect 7964 72176 7980 72240
rect 8044 72176 8060 72240
rect 8124 72176 8140 72240
rect 8204 72176 8220 72240
rect 8284 72236 13740 72240
rect 8284 72180 8375 72236
rect 8431 72180 11265 72236
rect 11321 72180 13740 72236
rect 8284 72176 13740 72180
rect 13804 72176 13820 72240
rect 13884 72176 13900 72240
rect 13964 72176 13980 72240
rect 14044 72176 14060 72240
rect 14124 72176 14140 72240
rect 14204 72236 14220 72240
rect 14211 72180 14220 72236
rect 14204 72176 14220 72180
rect 14284 72236 19740 72240
rect 14284 72180 17045 72236
rect 17101 72180 19740 72236
rect 14284 72176 19740 72180
rect 19804 72176 19820 72240
rect 19884 72176 19900 72240
rect 19964 72236 19980 72240
rect 19964 72176 19980 72180
rect 20044 72176 20060 72240
rect 20124 72176 20140 72240
rect 20204 72176 20220 72240
rect 20284 72236 25740 72240
rect 20284 72180 22825 72236
rect 22881 72180 25715 72236
rect 20284 72176 25740 72180
rect 25804 72176 25820 72240
rect 25884 72176 25900 72240
rect 25964 72176 25980 72240
rect 26044 72176 26060 72240
rect 26124 72176 26140 72240
rect 26204 72176 26220 72240
rect 26284 72236 31740 72240
rect 26284 72180 28605 72236
rect 28661 72180 31495 72236
rect 31551 72180 31740 72236
rect 26284 72176 31740 72180
rect 31804 72176 31820 72240
rect 31884 72176 31900 72240
rect 31964 72176 31980 72240
rect 32044 72176 32060 72240
rect 32124 72176 32140 72240
rect 32204 72176 32220 72240
rect 32284 72236 37740 72240
rect 32284 72180 34385 72236
rect 34441 72180 37275 72236
rect 37331 72180 37740 72236
rect 32284 72176 37740 72180
rect 37804 72176 37820 72240
rect 37884 72176 37900 72240
rect 37964 72176 37980 72240
rect 38044 72176 38060 72240
rect 38124 72176 38140 72240
rect 38204 72176 38220 72240
rect 38284 72236 43740 72240
rect 38284 72180 40165 72236
rect 40221 72180 43055 72236
rect 43111 72180 43740 72236
rect 38284 72176 43740 72180
rect 43804 72176 43820 72240
rect 43884 72176 43900 72240
rect 43964 72176 43980 72240
rect 44044 72176 44060 72240
rect 44124 72176 44140 72240
rect 44204 72176 44220 72240
rect 44284 72236 49740 72240
rect 49804 72236 49820 72240
rect 49884 72236 49900 72240
rect 44284 72180 45945 72236
rect 46001 72180 48892 72236
rect 48948 72180 49740 72236
rect 49810 72180 49820 72236
rect 49890 72180 49900 72236
rect 44284 72176 49740 72180
rect 49804 72176 49820 72180
rect 49884 72176 49900 72180
rect 49964 72176 49980 72240
rect 50044 72176 50060 72240
rect 50124 72176 50140 72240
rect 50204 72176 50220 72240
rect 50284 72236 55740 72240
rect 50284 72180 53048 72236
rect 53104 72180 53206 72236
rect 53262 72180 53562 72236
rect 53618 72180 54880 72236
rect 54936 72180 55473 72236
rect 55529 72180 55740 72236
rect 50284 72176 55740 72180
rect 55804 72176 55820 72240
rect 55884 72176 55900 72240
rect 55964 72176 55980 72240
rect 56044 72176 56060 72240
rect 56124 72176 56140 72240
rect 56204 72176 56220 72240
rect 56284 72236 61740 72240
rect 56284 72180 56619 72236
rect 56675 72180 58055 72236
rect 58111 72180 58135 72236
rect 58191 72180 59298 72236
rect 59354 72180 59456 72236
rect 59512 72180 59764 72236
rect 59820 72180 59910 72236
rect 59966 72180 60046 72236
rect 60102 72180 60126 72236
rect 60182 72180 61740 72236
rect 56284 72176 61740 72180
rect 61804 72176 61820 72240
rect 61884 72176 61900 72240
rect 61964 72176 61980 72240
rect 62044 72176 62060 72240
rect 62124 72176 62140 72240
rect 62204 72176 62220 72240
rect 62284 72236 67740 72240
rect 62284 72180 62418 72236
rect 62474 72180 62498 72236
rect 62554 72180 67740 72236
rect 62284 72176 67740 72180
rect 67804 72176 67820 72240
rect 67884 72176 67900 72240
rect 67964 72176 67980 72240
rect 68044 72176 68060 72240
rect 68124 72176 68140 72240
rect 68204 72176 68220 72240
rect 68284 72236 73740 72240
rect 68284 72180 71864 72236
rect 71920 72180 71944 72236
rect 72000 72180 72024 72236
rect 72080 72180 72104 72236
rect 72160 72180 73740 72236
rect 68284 72176 73740 72180
rect 73804 72176 73820 72240
rect 73884 72176 73900 72240
rect 73964 72176 73980 72240
rect 74044 72176 74060 72240
rect 74124 72176 74140 72240
rect 74204 72176 74220 72240
rect 74284 72176 75028 72240
rect 964 72160 75028 72176
rect 964 72096 1740 72160
rect 1804 72096 1820 72160
rect 1884 72096 1900 72160
rect 1964 72096 1980 72160
rect 2044 72096 2060 72160
rect 2124 72096 2140 72160
rect 2204 72096 2220 72160
rect 2284 72156 7740 72160
rect 2332 72100 2356 72156
rect 2412 72100 5485 72156
rect 5541 72100 7740 72156
rect 2284 72096 7740 72100
rect 7804 72096 7820 72160
rect 7884 72096 7900 72160
rect 7964 72096 7980 72160
rect 8044 72096 8060 72160
rect 8124 72096 8140 72160
rect 8204 72096 8220 72160
rect 8284 72156 13740 72160
rect 8284 72100 8375 72156
rect 8431 72100 11265 72156
rect 11321 72100 13740 72156
rect 8284 72096 13740 72100
rect 13804 72096 13820 72160
rect 13884 72096 13900 72160
rect 13964 72096 13980 72160
rect 14044 72096 14060 72160
rect 14124 72096 14140 72160
rect 14204 72156 14220 72160
rect 14211 72100 14220 72156
rect 14204 72096 14220 72100
rect 14284 72156 19740 72160
rect 14284 72100 17045 72156
rect 17101 72100 19740 72156
rect 14284 72096 19740 72100
rect 19804 72096 19820 72160
rect 19884 72096 19900 72160
rect 19964 72156 19980 72160
rect 19964 72096 19980 72100
rect 20044 72096 20060 72160
rect 20124 72096 20140 72160
rect 20204 72096 20220 72160
rect 20284 72156 25740 72160
rect 20284 72100 22825 72156
rect 22881 72100 25715 72156
rect 20284 72096 25740 72100
rect 25804 72096 25820 72160
rect 25884 72096 25900 72160
rect 25964 72096 25980 72160
rect 26044 72096 26060 72160
rect 26124 72096 26140 72160
rect 26204 72096 26220 72160
rect 26284 72156 31740 72160
rect 26284 72100 28605 72156
rect 28661 72100 31495 72156
rect 31551 72100 31740 72156
rect 26284 72096 31740 72100
rect 31804 72096 31820 72160
rect 31884 72096 31900 72160
rect 31964 72096 31980 72160
rect 32044 72096 32060 72160
rect 32124 72096 32140 72160
rect 32204 72096 32220 72160
rect 32284 72156 37740 72160
rect 32284 72100 34385 72156
rect 34441 72100 37275 72156
rect 37331 72100 37740 72156
rect 32284 72096 37740 72100
rect 37804 72096 37820 72160
rect 37884 72096 37900 72160
rect 37964 72096 37980 72160
rect 38044 72096 38060 72160
rect 38124 72096 38140 72160
rect 38204 72096 38220 72160
rect 38284 72156 43740 72160
rect 38284 72100 40165 72156
rect 40221 72100 43055 72156
rect 43111 72100 43740 72156
rect 38284 72096 43740 72100
rect 43804 72096 43820 72160
rect 43884 72096 43900 72160
rect 43964 72096 43980 72160
rect 44044 72096 44060 72160
rect 44124 72096 44140 72160
rect 44204 72096 44220 72160
rect 44284 72156 49740 72160
rect 49804 72156 49820 72160
rect 49884 72156 49900 72160
rect 44284 72100 45945 72156
rect 46001 72100 48892 72156
rect 48948 72100 49740 72156
rect 49810 72100 49820 72156
rect 49890 72100 49900 72156
rect 44284 72096 49740 72100
rect 49804 72096 49820 72100
rect 49884 72096 49900 72100
rect 49964 72096 49980 72160
rect 50044 72096 50060 72160
rect 50124 72096 50140 72160
rect 50204 72096 50220 72160
rect 50284 72156 55740 72160
rect 50284 72100 53048 72156
rect 53104 72100 53206 72156
rect 53262 72100 53562 72156
rect 53618 72100 54880 72156
rect 54936 72100 55473 72156
rect 55529 72100 55740 72156
rect 50284 72096 55740 72100
rect 55804 72096 55820 72160
rect 55884 72096 55900 72160
rect 55964 72096 55980 72160
rect 56044 72096 56060 72160
rect 56124 72096 56140 72160
rect 56204 72096 56220 72160
rect 56284 72156 61740 72160
rect 56284 72100 56619 72156
rect 56675 72100 58055 72156
rect 58111 72100 58135 72156
rect 58191 72100 59298 72156
rect 59354 72100 59456 72156
rect 59512 72100 59764 72156
rect 59820 72100 59910 72156
rect 59966 72100 60046 72156
rect 60102 72100 60126 72156
rect 60182 72100 61740 72156
rect 56284 72096 61740 72100
rect 61804 72096 61820 72160
rect 61884 72096 61900 72160
rect 61964 72096 61980 72160
rect 62044 72096 62060 72160
rect 62124 72096 62140 72160
rect 62204 72096 62220 72160
rect 62284 72156 67740 72160
rect 62284 72100 62418 72156
rect 62474 72100 62498 72156
rect 62554 72100 67740 72156
rect 62284 72096 67740 72100
rect 67804 72096 67820 72160
rect 67884 72096 67900 72160
rect 67964 72096 67980 72160
rect 68044 72096 68060 72160
rect 68124 72096 68140 72160
rect 68204 72096 68220 72160
rect 68284 72156 73740 72160
rect 68284 72100 71864 72156
rect 71920 72100 71944 72156
rect 72000 72100 72024 72156
rect 72080 72100 72104 72156
rect 72160 72100 73740 72156
rect 68284 72096 73740 72100
rect 73804 72096 73820 72160
rect 73884 72096 73900 72160
rect 73964 72096 73980 72160
rect 74044 72096 74060 72160
rect 74124 72096 74140 72160
rect 74204 72096 74220 72160
rect 74284 72096 75028 72160
rect 964 72080 75028 72096
rect 964 72016 1740 72080
rect 1804 72016 1820 72080
rect 1884 72016 1900 72080
rect 1964 72016 1980 72080
rect 2044 72016 2060 72080
rect 2124 72016 2140 72080
rect 2204 72016 2220 72080
rect 2284 72076 7740 72080
rect 2332 72020 2356 72076
rect 2412 72020 5485 72076
rect 5541 72020 7740 72076
rect 2284 72016 7740 72020
rect 7804 72016 7820 72080
rect 7884 72016 7900 72080
rect 7964 72016 7980 72080
rect 8044 72016 8060 72080
rect 8124 72016 8140 72080
rect 8204 72016 8220 72080
rect 8284 72076 13740 72080
rect 8284 72020 8375 72076
rect 8431 72020 11265 72076
rect 11321 72020 13740 72076
rect 8284 72016 13740 72020
rect 13804 72016 13820 72080
rect 13884 72016 13900 72080
rect 13964 72016 13980 72080
rect 14044 72016 14060 72080
rect 14124 72016 14140 72080
rect 14204 72076 14220 72080
rect 14211 72020 14220 72076
rect 14204 72016 14220 72020
rect 14284 72076 19740 72080
rect 14284 72020 17045 72076
rect 17101 72020 19740 72076
rect 14284 72016 19740 72020
rect 19804 72016 19820 72080
rect 19884 72016 19900 72080
rect 19964 72076 19980 72080
rect 19964 72016 19980 72020
rect 20044 72016 20060 72080
rect 20124 72016 20140 72080
rect 20204 72016 20220 72080
rect 20284 72076 25740 72080
rect 20284 72020 22825 72076
rect 22881 72020 25715 72076
rect 20284 72016 25740 72020
rect 25804 72016 25820 72080
rect 25884 72016 25900 72080
rect 25964 72016 25980 72080
rect 26044 72016 26060 72080
rect 26124 72016 26140 72080
rect 26204 72016 26220 72080
rect 26284 72076 31740 72080
rect 26284 72020 28605 72076
rect 28661 72020 31495 72076
rect 31551 72020 31740 72076
rect 26284 72016 31740 72020
rect 31804 72016 31820 72080
rect 31884 72016 31900 72080
rect 31964 72016 31980 72080
rect 32044 72016 32060 72080
rect 32124 72016 32140 72080
rect 32204 72016 32220 72080
rect 32284 72076 37740 72080
rect 32284 72020 34385 72076
rect 34441 72020 37275 72076
rect 37331 72020 37740 72076
rect 32284 72016 37740 72020
rect 37804 72016 37820 72080
rect 37884 72016 37900 72080
rect 37964 72016 37980 72080
rect 38044 72016 38060 72080
rect 38124 72016 38140 72080
rect 38204 72016 38220 72080
rect 38284 72076 43740 72080
rect 38284 72020 40165 72076
rect 40221 72020 43055 72076
rect 43111 72020 43740 72076
rect 38284 72016 43740 72020
rect 43804 72016 43820 72080
rect 43884 72016 43900 72080
rect 43964 72016 43980 72080
rect 44044 72016 44060 72080
rect 44124 72016 44140 72080
rect 44204 72016 44220 72080
rect 44284 72076 49740 72080
rect 49804 72076 49820 72080
rect 49884 72076 49900 72080
rect 44284 72020 45945 72076
rect 46001 72020 48892 72076
rect 48948 72020 49740 72076
rect 49810 72020 49820 72076
rect 49890 72020 49900 72076
rect 44284 72016 49740 72020
rect 49804 72016 49820 72020
rect 49884 72016 49900 72020
rect 49964 72016 49980 72080
rect 50044 72016 50060 72080
rect 50124 72016 50140 72080
rect 50204 72016 50220 72080
rect 50284 72076 55740 72080
rect 50284 72020 53048 72076
rect 53104 72020 53206 72076
rect 53262 72020 53562 72076
rect 53618 72020 54880 72076
rect 54936 72020 55473 72076
rect 55529 72020 55740 72076
rect 50284 72016 55740 72020
rect 55804 72016 55820 72080
rect 55884 72016 55900 72080
rect 55964 72016 55980 72080
rect 56044 72016 56060 72080
rect 56124 72016 56140 72080
rect 56204 72016 56220 72080
rect 56284 72076 61740 72080
rect 56284 72020 56619 72076
rect 56675 72020 58055 72076
rect 58111 72020 58135 72076
rect 58191 72020 59298 72076
rect 59354 72020 59456 72076
rect 59512 72020 59764 72076
rect 59820 72020 59910 72076
rect 59966 72020 60046 72076
rect 60102 72020 60126 72076
rect 60182 72020 61740 72076
rect 56284 72016 61740 72020
rect 61804 72016 61820 72080
rect 61884 72016 61900 72080
rect 61964 72016 61980 72080
rect 62044 72016 62060 72080
rect 62124 72016 62140 72080
rect 62204 72016 62220 72080
rect 62284 72076 67740 72080
rect 62284 72020 62418 72076
rect 62474 72020 62498 72076
rect 62554 72020 67740 72076
rect 62284 72016 67740 72020
rect 67804 72016 67820 72080
rect 67884 72016 67900 72080
rect 67964 72016 67980 72080
rect 68044 72016 68060 72080
rect 68124 72016 68140 72080
rect 68204 72016 68220 72080
rect 68284 72076 73740 72080
rect 68284 72020 71864 72076
rect 71920 72020 71944 72076
rect 72000 72020 72024 72076
rect 72080 72020 72104 72076
rect 72160 72020 73740 72076
rect 68284 72016 73740 72020
rect 73804 72016 73820 72080
rect 73884 72016 73900 72080
rect 73964 72016 73980 72080
rect 74044 72016 74060 72080
rect 74124 72016 74140 72080
rect 74204 72016 74220 72080
rect 74284 72016 75028 72080
rect 964 72000 75028 72016
rect 964 71936 1740 72000
rect 1804 71936 1820 72000
rect 1884 71936 1900 72000
rect 1964 71936 1980 72000
rect 2044 71936 2060 72000
rect 2124 71936 2140 72000
rect 2204 71936 2220 72000
rect 2284 71996 7740 72000
rect 2332 71940 2356 71996
rect 2412 71940 5485 71996
rect 5541 71940 7740 71996
rect 2284 71936 7740 71940
rect 7804 71936 7820 72000
rect 7884 71936 7900 72000
rect 7964 71936 7980 72000
rect 8044 71936 8060 72000
rect 8124 71936 8140 72000
rect 8204 71936 8220 72000
rect 8284 71996 13740 72000
rect 8284 71940 8375 71996
rect 8431 71940 11265 71996
rect 11321 71940 13740 71996
rect 8284 71936 13740 71940
rect 13804 71936 13820 72000
rect 13884 71936 13900 72000
rect 13964 71936 13980 72000
rect 14044 71936 14060 72000
rect 14124 71936 14140 72000
rect 14204 71996 14220 72000
rect 14211 71940 14220 71996
rect 14204 71936 14220 71940
rect 14284 71996 19740 72000
rect 14284 71940 17045 71996
rect 17101 71940 19740 71996
rect 14284 71936 19740 71940
rect 19804 71936 19820 72000
rect 19884 71936 19900 72000
rect 19964 71996 19980 72000
rect 19964 71936 19980 71940
rect 20044 71936 20060 72000
rect 20124 71936 20140 72000
rect 20204 71936 20220 72000
rect 20284 71996 25740 72000
rect 20284 71940 22825 71996
rect 22881 71940 25715 71996
rect 20284 71936 25740 71940
rect 25804 71936 25820 72000
rect 25884 71936 25900 72000
rect 25964 71936 25980 72000
rect 26044 71936 26060 72000
rect 26124 71936 26140 72000
rect 26204 71936 26220 72000
rect 26284 71996 31740 72000
rect 26284 71940 28605 71996
rect 28661 71940 31495 71996
rect 31551 71940 31740 71996
rect 26284 71936 31740 71940
rect 31804 71936 31820 72000
rect 31884 71936 31900 72000
rect 31964 71936 31980 72000
rect 32044 71936 32060 72000
rect 32124 71936 32140 72000
rect 32204 71936 32220 72000
rect 32284 71996 37740 72000
rect 32284 71940 34385 71996
rect 34441 71940 37275 71996
rect 37331 71940 37740 71996
rect 32284 71936 37740 71940
rect 37804 71936 37820 72000
rect 37884 71936 37900 72000
rect 37964 71936 37980 72000
rect 38044 71936 38060 72000
rect 38124 71936 38140 72000
rect 38204 71936 38220 72000
rect 38284 71996 43740 72000
rect 38284 71940 40165 71996
rect 40221 71940 43055 71996
rect 43111 71940 43740 71996
rect 38284 71936 43740 71940
rect 43804 71936 43820 72000
rect 43884 71936 43900 72000
rect 43964 71936 43980 72000
rect 44044 71936 44060 72000
rect 44124 71936 44140 72000
rect 44204 71936 44220 72000
rect 44284 71996 49740 72000
rect 49804 71996 49820 72000
rect 49884 71996 49900 72000
rect 44284 71940 45945 71996
rect 46001 71940 48892 71996
rect 48948 71940 49740 71996
rect 49810 71940 49820 71996
rect 49890 71940 49900 71996
rect 44284 71936 49740 71940
rect 49804 71936 49820 71940
rect 49884 71936 49900 71940
rect 49964 71936 49980 72000
rect 50044 71936 50060 72000
rect 50124 71936 50140 72000
rect 50204 71936 50220 72000
rect 50284 71996 55740 72000
rect 50284 71940 53048 71996
rect 53104 71940 53206 71996
rect 53262 71940 53562 71996
rect 53618 71940 54880 71996
rect 54936 71940 55473 71996
rect 55529 71940 55740 71996
rect 50284 71936 55740 71940
rect 55804 71936 55820 72000
rect 55884 71936 55900 72000
rect 55964 71936 55980 72000
rect 56044 71936 56060 72000
rect 56124 71936 56140 72000
rect 56204 71936 56220 72000
rect 56284 71996 61740 72000
rect 56284 71940 56619 71996
rect 56675 71940 58055 71996
rect 58111 71940 58135 71996
rect 58191 71940 59298 71996
rect 59354 71940 59456 71996
rect 59512 71940 59764 71996
rect 59820 71940 59910 71996
rect 59966 71940 60046 71996
rect 60102 71940 60126 71996
rect 60182 71940 61740 71996
rect 56284 71936 61740 71940
rect 61804 71936 61820 72000
rect 61884 71936 61900 72000
rect 61964 71936 61980 72000
rect 62044 71936 62060 72000
rect 62124 71936 62140 72000
rect 62204 71936 62220 72000
rect 62284 71996 67740 72000
rect 62284 71940 62418 71996
rect 62474 71940 62498 71996
rect 62554 71940 67740 71996
rect 62284 71936 67740 71940
rect 67804 71936 67820 72000
rect 67884 71936 67900 72000
rect 67964 71936 67980 72000
rect 68044 71936 68060 72000
rect 68124 71936 68140 72000
rect 68204 71936 68220 72000
rect 68284 71996 73740 72000
rect 68284 71940 71864 71996
rect 71920 71940 71944 71996
rect 72000 71940 72024 71996
rect 72080 71940 72104 71996
rect 72160 71940 73740 71996
rect 68284 71936 73740 71940
rect 73804 71936 73820 72000
rect 73884 71936 73900 72000
rect 73964 71936 73980 72000
rect 74044 71936 74060 72000
rect 74124 71936 74140 72000
rect 74204 71936 74220 72000
rect 74284 71936 75028 72000
rect 964 71912 75028 71936
rect 63493 65244 63559 65245
rect 63493 65242 63540 65244
rect 63448 65240 63540 65242
rect 63448 65184 63498 65240
rect 63448 65182 63540 65184
rect 63493 65180 63540 65182
rect 63604 65180 63610 65244
rect 63493 65179 63559 65180
rect 964 64592 75028 64616
rect 964 64588 4740 64592
rect 964 64532 2136 64588
rect 2192 64532 4740 64588
rect 964 64528 4740 64532
rect 4804 64528 4820 64592
rect 4884 64528 4900 64592
rect 4964 64528 4980 64592
rect 5044 64528 5060 64592
rect 5124 64528 5140 64592
rect 5204 64528 5220 64592
rect 5284 64588 10740 64592
rect 5284 64532 5632 64588
rect 5688 64532 8522 64588
rect 8578 64532 10740 64588
rect 5284 64528 10740 64532
rect 10804 64528 10820 64592
rect 10884 64528 10900 64592
rect 10964 64528 10980 64592
rect 11044 64528 11060 64592
rect 11124 64528 11140 64592
rect 11204 64528 11220 64592
rect 11284 64588 16740 64592
rect 11284 64532 11412 64588
rect 11468 64532 14302 64588
rect 14358 64532 16740 64588
rect 11284 64528 16740 64532
rect 16804 64528 16820 64592
rect 16884 64528 16900 64592
rect 16964 64528 16980 64592
rect 17044 64528 17060 64592
rect 17124 64528 17140 64592
rect 17204 64588 17220 64592
rect 17284 64588 22740 64592
rect 17284 64532 20082 64588
rect 20138 64532 22740 64588
rect 17204 64528 17220 64532
rect 17284 64528 22740 64532
rect 22804 64528 22820 64592
rect 22884 64528 22900 64592
rect 22964 64588 22980 64592
rect 22964 64532 22972 64588
rect 22964 64528 22980 64532
rect 23044 64528 23060 64592
rect 23124 64528 23140 64592
rect 23204 64528 23220 64592
rect 23284 64588 28740 64592
rect 28804 64588 28820 64592
rect 23284 64532 25862 64588
rect 25918 64532 28740 64588
rect 28808 64532 28820 64588
rect 23284 64528 28740 64532
rect 28804 64528 28820 64532
rect 28884 64528 28900 64592
rect 28964 64528 28980 64592
rect 29044 64528 29060 64592
rect 29124 64528 29140 64592
rect 29204 64528 29220 64592
rect 29284 64588 34740 64592
rect 29284 64532 31642 64588
rect 31698 64532 34532 64588
rect 34588 64532 34740 64588
rect 29284 64528 34740 64532
rect 34804 64528 34820 64592
rect 34884 64528 34900 64592
rect 34964 64528 34980 64592
rect 35044 64528 35060 64592
rect 35124 64528 35140 64592
rect 35204 64528 35220 64592
rect 35284 64588 40740 64592
rect 35284 64532 37422 64588
rect 37478 64532 40312 64588
rect 40368 64532 40740 64588
rect 35284 64528 40740 64532
rect 40804 64528 40820 64592
rect 40884 64528 40900 64592
rect 40964 64528 40980 64592
rect 41044 64528 41060 64592
rect 41124 64528 41140 64592
rect 41204 64528 41220 64592
rect 41284 64588 46740 64592
rect 41284 64532 43202 64588
rect 43258 64532 46092 64588
rect 46148 64532 46740 64588
rect 41284 64528 46740 64532
rect 46804 64528 46820 64592
rect 46884 64528 46900 64592
rect 46964 64528 46980 64592
rect 47044 64528 47060 64592
rect 47124 64528 47140 64592
rect 47204 64528 47220 64592
rect 47284 64588 52740 64592
rect 47284 64532 49100 64588
rect 49156 64532 52329 64588
rect 52385 64532 52740 64588
rect 47284 64528 52740 64532
rect 52804 64528 52820 64592
rect 52884 64528 52900 64592
rect 52964 64528 52980 64592
rect 53044 64528 53060 64592
rect 53124 64528 53140 64592
rect 53204 64528 53220 64592
rect 53284 64588 58740 64592
rect 53284 64532 53730 64588
rect 53786 64532 53898 64588
rect 53954 64532 54642 64588
rect 54698 64532 55032 64588
rect 55088 64532 55748 64588
rect 55804 64532 56326 64588
rect 56382 64532 56771 64588
rect 56827 64532 57075 64588
rect 57131 64532 57917 64588
rect 57973 64532 58557 64588
rect 58613 64532 58740 64588
rect 53284 64528 58740 64532
rect 58804 64528 58820 64592
rect 58884 64528 58900 64592
rect 58964 64528 58980 64592
rect 59044 64528 59060 64592
rect 59124 64528 59140 64592
rect 59204 64528 59220 64592
rect 59284 64588 64740 64592
rect 59284 64532 60418 64588
rect 60474 64532 60576 64588
rect 60632 64532 62620 64588
rect 62676 64532 62700 64588
rect 62756 64532 64740 64588
rect 59284 64528 64740 64532
rect 64804 64528 64820 64592
rect 64884 64528 64900 64592
rect 64964 64528 64980 64592
rect 65044 64528 65060 64592
rect 65124 64528 65140 64592
rect 65204 64528 65220 64592
rect 65284 64528 70740 64592
rect 70804 64528 70820 64592
rect 70884 64528 70900 64592
rect 70964 64528 70980 64592
rect 71044 64528 71060 64592
rect 71124 64528 71140 64592
rect 71204 64528 71220 64592
rect 71284 64588 75028 64592
rect 71284 64532 74216 64588
rect 74272 64532 74296 64588
rect 74352 64532 74376 64588
rect 74432 64532 74456 64588
rect 74512 64532 75028 64588
rect 71284 64528 75028 64532
rect 964 64512 75028 64528
rect 964 64508 4740 64512
rect 964 64452 2136 64508
rect 2192 64452 4740 64508
rect 964 64448 4740 64452
rect 4804 64448 4820 64512
rect 4884 64448 4900 64512
rect 4964 64448 4980 64512
rect 5044 64448 5060 64512
rect 5124 64448 5140 64512
rect 5204 64448 5220 64512
rect 5284 64508 10740 64512
rect 5284 64452 5632 64508
rect 5688 64452 8522 64508
rect 8578 64452 10740 64508
rect 5284 64448 10740 64452
rect 10804 64448 10820 64512
rect 10884 64448 10900 64512
rect 10964 64448 10980 64512
rect 11044 64448 11060 64512
rect 11124 64448 11140 64512
rect 11204 64448 11220 64512
rect 11284 64508 16740 64512
rect 11284 64452 11412 64508
rect 11468 64452 14302 64508
rect 14358 64452 16740 64508
rect 11284 64448 16740 64452
rect 16804 64448 16820 64512
rect 16884 64448 16900 64512
rect 16964 64448 16980 64512
rect 17044 64448 17060 64512
rect 17124 64448 17140 64512
rect 17204 64508 17220 64512
rect 17284 64508 22740 64512
rect 17284 64452 20082 64508
rect 20138 64452 22740 64508
rect 17204 64448 17220 64452
rect 17284 64448 22740 64452
rect 22804 64448 22820 64512
rect 22884 64448 22900 64512
rect 22964 64508 22980 64512
rect 22964 64452 22972 64508
rect 22964 64448 22980 64452
rect 23044 64448 23060 64512
rect 23124 64448 23140 64512
rect 23204 64448 23220 64512
rect 23284 64508 28740 64512
rect 28804 64508 28820 64512
rect 23284 64452 25862 64508
rect 25918 64452 28740 64508
rect 28808 64452 28820 64508
rect 23284 64448 28740 64452
rect 28804 64448 28820 64452
rect 28884 64448 28900 64512
rect 28964 64448 28980 64512
rect 29044 64448 29060 64512
rect 29124 64448 29140 64512
rect 29204 64448 29220 64512
rect 29284 64508 34740 64512
rect 29284 64452 31642 64508
rect 31698 64452 34532 64508
rect 34588 64452 34740 64508
rect 29284 64448 34740 64452
rect 34804 64448 34820 64512
rect 34884 64448 34900 64512
rect 34964 64448 34980 64512
rect 35044 64448 35060 64512
rect 35124 64448 35140 64512
rect 35204 64448 35220 64512
rect 35284 64508 40740 64512
rect 35284 64452 37422 64508
rect 37478 64452 40312 64508
rect 40368 64452 40740 64508
rect 35284 64448 40740 64452
rect 40804 64448 40820 64512
rect 40884 64448 40900 64512
rect 40964 64448 40980 64512
rect 41044 64448 41060 64512
rect 41124 64448 41140 64512
rect 41204 64448 41220 64512
rect 41284 64508 46740 64512
rect 41284 64452 43202 64508
rect 43258 64452 46092 64508
rect 46148 64452 46740 64508
rect 41284 64448 46740 64452
rect 46804 64448 46820 64512
rect 46884 64448 46900 64512
rect 46964 64448 46980 64512
rect 47044 64448 47060 64512
rect 47124 64448 47140 64512
rect 47204 64448 47220 64512
rect 47284 64508 52740 64512
rect 47284 64452 49100 64508
rect 49156 64452 52329 64508
rect 52385 64452 52740 64508
rect 47284 64448 52740 64452
rect 52804 64448 52820 64512
rect 52884 64448 52900 64512
rect 52964 64448 52980 64512
rect 53044 64448 53060 64512
rect 53124 64448 53140 64512
rect 53204 64448 53220 64512
rect 53284 64508 58740 64512
rect 53284 64452 53730 64508
rect 53786 64452 53898 64508
rect 53954 64452 54642 64508
rect 54698 64452 55032 64508
rect 55088 64452 55748 64508
rect 55804 64452 56326 64508
rect 56382 64452 56771 64508
rect 56827 64452 57075 64508
rect 57131 64452 57917 64508
rect 57973 64452 58557 64508
rect 58613 64452 58740 64508
rect 53284 64448 58740 64452
rect 58804 64448 58820 64512
rect 58884 64448 58900 64512
rect 58964 64448 58980 64512
rect 59044 64448 59060 64512
rect 59124 64448 59140 64512
rect 59204 64448 59220 64512
rect 59284 64508 64740 64512
rect 59284 64452 60418 64508
rect 60474 64452 60576 64508
rect 60632 64452 62620 64508
rect 62676 64452 62700 64508
rect 62756 64452 64740 64508
rect 59284 64448 64740 64452
rect 64804 64448 64820 64512
rect 64884 64448 64900 64512
rect 64964 64448 64980 64512
rect 65044 64448 65060 64512
rect 65124 64448 65140 64512
rect 65204 64448 65220 64512
rect 65284 64448 70740 64512
rect 70804 64448 70820 64512
rect 70884 64448 70900 64512
rect 70964 64448 70980 64512
rect 71044 64448 71060 64512
rect 71124 64448 71140 64512
rect 71204 64448 71220 64512
rect 71284 64508 75028 64512
rect 71284 64452 74216 64508
rect 74272 64452 74296 64508
rect 74352 64452 74376 64508
rect 74432 64452 74456 64508
rect 74512 64452 75028 64508
rect 71284 64448 75028 64452
rect 964 64432 75028 64448
rect 964 64428 4740 64432
rect 964 64372 2136 64428
rect 2192 64372 4740 64428
rect 964 64368 4740 64372
rect 4804 64368 4820 64432
rect 4884 64368 4900 64432
rect 4964 64368 4980 64432
rect 5044 64368 5060 64432
rect 5124 64368 5140 64432
rect 5204 64368 5220 64432
rect 5284 64428 10740 64432
rect 5284 64372 5632 64428
rect 5688 64372 8522 64428
rect 8578 64372 10740 64428
rect 5284 64368 10740 64372
rect 10804 64368 10820 64432
rect 10884 64368 10900 64432
rect 10964 64368 10980 64432
rect 11044 64368 11060 64432
rect 11124 64368 11140 64432
rect 11204 64368 11220 64432
rect 11284 64428 16740 64432
rect 11284 64372 11412 64428
rect 11468 64372 14302 64428
rect 14358 64372 16740 64428
rect 11284 64368 16740 64372
rect 16804 64368 16820 64432
rect 16884 64368 16900 64432
rect 16964 64368 16980 64432
rect 17044 64368 17060 64432
rect 17124 64368 17140 64432
rect 17204 64428 17220 64432
rect 17284 64428 22740 64432
rect 17284 64372 20082 64428
rect 20138 64372 22740 64428
rect 17204 64368 17220 64372
rect 17284 64368 22740 64372
rect 22804 64368 22820 64432
rect 22884 64368 22900 64432
rect 22964 64428 22980 64432
rect 22964 64372 22972 64428
rect 22964 64368 22980 64372
rect 23044 64368 23060 64432
rect 23124 64368 23140 64432
rect 23204 64368 23220 64432
rect 23284 64428 28740 64432
rect 28804 64428 28820 64432
rect 23284 64372 25862 64428
rect 25918 64372 28740 64428
rect 28808 64372 28820 64428
rect 23284 64368 28740 64372
rect 28804 64368 28820 64372
rect 28884 64368 28900 64432
rect 28964 64368 28980 64432
rect 29044 64368 29060 64432
rect 29124 64368 29140 64432
rect 29204 64368 29220 64432
rect 29284 64428 34740 64432
rect 29284 64372 31642 64428
rect 31698 64372 34532 64428
rect 34588 64372 34740 64428
rect 29284 64368 34740 64372
rect 34804 64368 34820 64432
rect 34884 64368 34900 64432
rect 34964 64368 34980 64432
rect 35044 64368 35060 64432
rect 35124 64368 35140 64432
rect 35204 64368 35220 64432
rect 35284 64428 40740 64432
rect 35284 64372 37422 64428
rect 37478 64372 40312 64428
rect 40368 64372 40740 64428
rect 35284 64368 40740 64372
rect 40804 64368 40820 64432
rect 40884 64368 40900 64432
rect 40964 64368 40980 64432
rect 41044 64368 41060 64432
rect 41124 64368 41140 64432
rect 41204 64368 41220 64432
rect 41284 64428 46740 64432
rect 41284 64372 43202 64428
rect 43258 64372 46092 64428
rect 46148 64372 46740 64428
rect 41284 64368 46740 64372
rect 46804 64368 46820 64432
rect 46884 64368 46900 64432
rect 46964 64368 46980 64432
rect 47044 64368 47060 64432
rect 47124 64368 47140 64432
rect 47204 64368 47220 64432
rect 47284 64428 52740 64432
rect 47284 64372 49100 64428
rect 49156 64372 52329 64428
rect 52385 64372 52740 64428
rect 47284 64368 52740 64372
rect 52804 64368 52820 64432
rect 52884 64368 52900 64432
rect 52964 64368 52980 64432
rect 53044 64368 53060 64432
rect 53124 64368 53140 64432
rect 53204 64368 53220 64432
rect 53284 64428 58740 64432
rect 53284 64372 53730 64428
rect 53786 64372 53898 64428
rect 53954 64372 54642 64428
rect 54698 64372 55032 64428
rect 55088 64372 55748 64428
rect 55804 64372 56326 64428
rect 56382 64372 56771 64428
rect 56827 64372 57075 64428
rect 57131 64372 57917 64428
rect 57973 64372 58557 64428
rect 58613 64372 58740 64428
rect 53284 64368 58740 64372
rect 58804 64368 58820 64432
rect 58884 64368 58900 64432
rect 58964 64368 58980 64432
rect 59044 64368 59060 64432
rect 59124 64368 59140 64432
rect 59204 64368 59220 64432
rect 59284 64428 64740 64432
rect 59284 64372 60418 64428
rect 60474 64372 60576 64428
rect 60632 64372 62620 64428
rect 62676 64372 62700 64428
rect 62756 64372 64740 64428
rect 59284 64368 64740 64372
rect 64804 64368 64820 64432
rect 64884 64368 64900 64432
rect 64964 64368 64980 64432
rect 65044 64368 65060 64432
rect 65124 64368 65140 64432
rect 65204 64368 65220 64432
rect 65284 64368 70740 64432
rect 70804 64368 70820 64432
rect 70884 64368 70900 64432
rect 70964 64368 70980 64432
rect 71044 64368 71060 64432
rect 71124 64368 71140 64432
rect 71204 64368 71220 64432
rect 71284 64428 75028 64432
rect 71284 64372 74216 64428
rect 74272 64372 74296 64428
rect 74352 64372 74376 64428
rect 74432 64372 74456 64428
rect 74512 64372 75028 64428
rect 71284 64368 75028 64372
rect 964 64352 75028 64368
rect 964 64348 4740 64352
rect 964 64292 2136 64348
rect 2192 64292 4740 64348
rect 964 64288 4740 64292
rect 4804 64288 4820 64352
rect 4884 64288 4900 64352
rect 4964 64288 4980 64352
rect 5044 64288 5060 64352
rect 5124 64288 5140 64352
rect 5204 64288 5220 64352
rect 5284 64348 10740 64352
rect 5284 64292 5632 64348
rect 5688 64292 8522 64348
rect 8578 64292 10740 64348
rect 5284 64288 10740 64292
rect 10804 64288 10820 64352
rect 10884 64288 10900 64352
rect 10964 64288 10980 64352
rect 11044 64288 11060 64352
rect 11124 64288 11140 64352
rect 11204 64288 11220 64352
rect 11284 64348 16740 64352
rect 11284 64292 11412 64348
rect 11468 64292 14302 64348
rect 14358 64292 16740 64348
rect 11284 64288 16740 64292
rect 16804 64288 16820 64352
rect 16884 64288 16900 64352
rect 16964 64288 16980 64352
rect 17044 64288 17060 64352
rect 17124 64288 17140 64352
rect 17204 64348 17220 64352
rect 17284 64348 22740 64352
rect 17284 64292 20082 64348
rect 20138 64292 22740 64348
rect 17204 64288 17220 64292
rect 17284 64288 22740 64292
rect 22804 64288 22820 64352
rect 22884 64288 22900 64352
rect 22964 64348 22980 64352
rect 22964 64292 22972 64348
rect 22964 64288 22980 64292
rect 23044 64288 23060 64352
rect 23124 64288 23140 64352
rect 23204 64288 23220 64352
rect 23284 64348 28740 64352
rect 28804 64348 28820 64352
rect 23284 64292 25862 64348
rect 25918 64292 28740 64348
rect 28808 64292 28820 64348
rect 23284 64288 28740 64292
rect 28804 64288 28820 64292
rect 28884 64288 28900 64352
rect 28964 64288 28980 64352
rect 29044 64288 29060 64352
rect 29124 64288 29140 64352
rect 29204 64288 29220 64352
rect 29284 64348 34740 64352
rect 29284 64292 31642 64348
rect 31698 64292 34532 64348
rect 34588 64292 34740 64348
rect 29284 64288 34740 64292
rect 34804 64288 34820 64352
rect 34884 64288 34900 64352
rect 34964 64288 34980 64352
rect 35044 64288 35060 64352
rect 35124 64288 35140 64352
rect 35204 64288 35220 64352
rect 35284 64348 40740 64352
rect 35284 64292 37422 64348
rect 37478 64292 40312 64348
rect 40368 64292 40740 64348
rect 35284 64288 40740 64292
rect 40804 64288 40820 64352
rect 40884 64288 40900 64352
rect 40964 64288 40980 64352
rect 41044 64288 41060 64352
rect 41124 64288 41140 64352
rect 41204 64288 41220 64352
rect 41284 64348 46740 64352
rect 41284 64292 43202 64348
rect 43258 64292 46092 64348
rect 46148 64292 46740 64348
rect 41284 64288 46740 64292
rect 46804 64288 46820 64352
rect 46884 64288 46900 64352
rect 46964 64288 46980 64352
rect 47044 64288 47060 64352
rect 47124 64288 47140 64352
rect 47204 64288 47220 64352
rect 47284 64348 52740 64352
rect 47284 64292 49100 64348
rect 49156 64292 52329 64348
rect 52385 64292 52740 64348
rect 47284 64288 52740 64292
rect 52804 64288 52820 64352
rect 52884 64288 52900 64352
rect 52964 64288 52980 64352
rect 53044 64288 53060 64352
rect 53124 64288 53140 64352
rect 53204 64288 53220 64352
rect 53284 64348 58740 64352
rect 53284 64292 53730 64348
rect 53786 64292 53898 64348
rect 53954 64292 54642 64348
rect 54698 64292 55032 64348
rect 55088 64292 55748 64348
rect 55804 64292 56326 64348
rect 56382 64292 56771 64348
rect 56827 64292 57075 64348
rect 57131 64292 57917 64348
rect 57973 64292 58557 64348
rect 58613 64292 58740 64348
rect 53284 64288 58740 64292
rect 58804 64288 58820 64352
rect 58884 64288 58900 64352
rect 58964 64288 58980 64352
rect 59044 64288 59060 64352
rect 59124 64288 59140 64352
rect 59204 64288 59220 64352
rect 59284 64348 64740 64352
rect 59284 64292 60418 64348
rect 60474 64292 60576 64348
rect 60632 64292 62620 64348
rect 62676 64292 62700 64348
rect 62756 64292 64740 64348
rect 59284 64288 64740 64292
rect 64804 64288 64820 64352
rect 64884 64288 64900 64352
rect 64964 64288 64980 64352
rect 65044 64288 65060 64352
rect 65124 64288 65140 64352
rect 65204 64288 65220 64352
rect 65284 64288 70740 64352
rect 70804 64288 70820 64352
rect 70884 64288 70900 64352
rect 70964 64288 70980 64352
rect 71044 64288 71060 64352
rect 71124 64288 71140 64352
rect 71204 64288 71220 64352
rect 71284 64348 75028 64352
rect 71284 64292 74216 64348
rect 74272 64292 74296 64348
rect 74352 64292 74376 64348
rect 74432 64292 74456 64348
rect 74512 64292 75028 64348
rect 71284 64288 75028 64292
rect 964 64264 75028 64288
rect 63493 63202 63559 63205
rect 63718 63202 63724 63204
rect 63493 63200 63724 63202
rect 63493 63144 63498 63200
rect 63554 63144 63724 63200
rect 63493 63142 63724 63144
rect 63493 63139 63559 63142
rect 63718 63140 63724 63142
rect 63788 63140 63794 63204
rect 964 62240 75028 62264
rect 964 62176 1740 62240
rect 1804 62176 1820 62240
rect 1884 62176 1900 62240
rect 1964 62176 1980 62240
rect 2044 62176 2060 62240
rect 2124 62176 2140 62240
rect 2204 62176 2220 62240
rect 2284 62236 7740 62240
rect 2332 62180 2356 62236
rect 2412 62180 5485 62236
rect 5541 62180 7740 62236
rect 2284 62176 7740 62180
rect 7804 62176 7820 62240
rect 7884 62176 7900 62240
rect 7964 62176 7980 62240
rect 8044 62176 8060 62240
rect 8124 62176 8140 62240
rect 8204 62176 8220 62240
rect 8284 62236 13740 62240
rect 8284 62180 8375 62236
rect 8431 62180 11265 62236
rect 11321 62180 13740 62236
rect 8284 62176 13740 62180
rect 13804 62176 13820 62240
rect 13884 62176 13900 62240
rect 13964 62176 13980 62240
rect 14044 62176 14060 62240
rect 14124 62176 14140 62240
rect 14204 62236 14220 62240
rect 14211 62180 14220 62236
rect 14204 62176 14220 62180
rect 14284 62236 19740 62240
rect 14284 62180 17045 62236
rect 17101 62180 19740 62236
rect 14284 62176 19740 62180
rect 19804 62176 19820 62240
rect 19884 62176 19900 62240
rect 19964 62236 19980 62240
rect 19964 62176 19980 62180
rect 20044 62176 20060 62240
rect 20124 62176 20140 62240
rect 20204 62176 20220 62240
rect 20284 62236 25740 62240
rect 20284 62180 22825 62236
rect 22881 62180 25715 62236
rect 20284 62176 25740 62180
rect 25804 62176 25820 62240
rect 25884 62176 25900 62240
rect 25964 62176 25980 62240
rect 26044 62176 26060 62240
rect 26124 62176 26140 62240
rect 26204 62176 26220 62240
rect 26284 62236 31740 62240
rect 26284 62180 28605 62236
rect 28661 62180 31495 62236
rect 31551 62180 31740 62236
rect 26284 62176 31740 62180
rect 31804 62176 31820 62240
rect 31884 62176 31900 62240
rect 31964 62176 31980 62240
rect 32044 62176 32060 62240
rect 32124 62176 32140 62240
rect 32204 62176 32220 62240
rect 32284 62236 37740 62240
rect 32284 62180 34385 62236
rect 34441 62180 37275 62236
rect 37331 62180 37740 62236
rect 32284 62176 37740 62180
rect 37804 62176 37820 62240
rect 37884 62176 37900 62240
rect 37964 62176 37980 62240
rect 38044 62176 38060 62240
rect 38124 62176 38140 62240
rect 38204 62176 38220 62240
rect 38284 62236 43740 62240
rect 38284 62180 40165 62236
rect 40221 62180 43055 62236
rect 43111 62180 43740 62236
rect 38284 62176 43740 62180
rect 43804 62176 43820 62240
rect 43884 62176 43900 62240
rect 43964 62176 43980 62240
rect 44044 62176 44060 62240
rect 44124 62176 44140 62240
rect 44204 62176 44220 62240
rect 44284 62236 49740 62240
rect 49804 62236 49820 62240
rect 49884 62236 49900 62240
rect 44284 62180 45945 62236
rect 46001 62180 48892 62236
rect 48948 62180 49740 62236
rect 49810 62180 49820 62236
rect 49890 62180 49900 62236
rect 44284 62176 49740 62180
rect 49804 62176 49820 62180
rect 49884 62176 49900 62180
rect 49964 62176 49980 62240
rect 50044 62176 50060 62240
rect 50124 62176 50140 62240
rect 50204 62176 50220 62240
rect 50284 62236 55740 62240
rect 50284 62180 53048 62236
rect 53104 62180 53206 62236
rect 53262 62180 53562 62236
rect 53618 62180 54880 62236
rect 54936 62180 55473 62236
rect 55529 62180 55740 62236
rect 50284 62176 55740 62180
rect 55804 62176 55820 62240
rect 55884 62176 55900 62240
rect 55964 62176 55980 62240
rect 56044 62176 56060 62240
rect 56124 62176 56140 62240
rect 56204 62176 56220 62240
rect 56284 62236 61740 62240
rect 56284 62180 56619 62236
rect 56675 62180 58055 62236
rect 58111 62180 58135 62236
rect 58191 62180 59298 62236
rect 59354 62180 59456 62236
rect 59512 62180 59764 62236
rect 59820 62180 59910 62236
rect 59966 62180 60046 62236
rect 60102 62180 60126 62236
rect 60182 62180 61740 62236
rect 56284 62176 61740 62180
rect 61804 62176 61820 62240
rect 61884 62176 61900 62240
rect 61964 62176 61980 62240
rect 62044 62176 62060 62240
rect 62124 62176 62140 62240
rect 62204 62176 62220 62240
rect 62284 62236 67740 62240
rect 62284 62180 62418 62236
rect 62474 62180 62498 62236
rect 62554 62180 67740 62236
rect 62284 62176 67740 62180
rect 67804 62176 67820 62240
rect 67884 62176 67900 62240
rect 67964 62176 67980 62240
rect 68044 62176 68060 62240
rect 68124 62176 68140 62240
rect 68204 62176 68220 62240
rect 68284 62236 73740 62240
rect 68284 62180 71864 62236
rect 71920 62180 71944 62236
rect 72000 62180 72024 62236
rect 72080 62180 72104 62236
rect 72160 62180 73740 62236
rect 68284 62176 73740 62180
rect 73804 62176 73820 62240
rect 73884 62176 73900 62240
rect 73964 62176 73980 62240
rect 74044 62176 74060 62240
rect 74124 62176 74140 62240
rect 74204 62176 74220 62240
rect 74284 62176 75028 62240
rect 964 62160 75028 62176
rect 964 62096 1740 62160
rect 1804 62096 1820 62160
rect 1884 62096 1900 62160
rect 1964 62096 1980 62160
rect 2044 62096 2060 62160
rect 2124 62096 2140 62160
rect 2204 62096 2220 62160
rect 2284 62156 7740 62160
rect 2332 62100 2356 62156
rect 2412 62100 5485 62156
rect 5541 62100 7740 62156
rect 2284 62096 7740 62100
rect 7804 62096 7820 62160
rect 7884 62096 7900 62160
rect 7964 62096 7980 62160
rect 8044 62096 8060 62160
rect 8124 62096 8140 62160
rect 8204 62096 8220 62160
rect 8284 62156 13740 62160
rect 8284 62100 8375 62156
rect 8431 62100 11265 62156
rect 11321 62100 13740 62156
rect 8284 62096 13740 62100
rect 13804 62096 13820 62160
rect 13884 62096 13900 62160
rect 13964 62096 13980 62160
rect 14044 62096 14060 62160
rect 14124 62096 14140 62160
rect 14204 62156 14220 62160
rect 14211 62100 14220 62156
rect 14204 62096 14220 62100
rect 14284 62156 19740 62160
rect 14284 62100 17045 62156
rect 17101 62100 19740 62156
rect 14284 62096 19740 62100
rect 19804 62096 19820 62160
rect 19884 62096 19900 62160
rect 19964 62156 19980 62160
rect 19964 62096 19980 62100
rect 20044 62096 20060 62160
rect 20124 62096 20140 62160
rect 20204 62096 20220 62160
rect 20284 62156 25740 62160
rect 20284 62100 22825 62156
rect 22881 62100 25715 62156
rect 20284 62096 25740 62100
rect 25804 62096 25820 62160
rect 25884 62096 25900 62160
rect 25964 62096 25980 62160
rect 26044 62096 26060 62160
rect 26124 62096 26140 62160
rect 26204 62096 26220 62160
rect 26284 62156 31740 62160
rect 26284 62100 28605 62156
rect 28661 62100 31495 62156
rect 31551 62100 31740 62156
rect 26284 62096 31740 62100
rect 31804 62096 31820 62160
rect 31884 62096 31900 62160
rect 31964 62096 31980 62160
rect 32044 62096 32060 62160
rect 32124 62096 32140 62160
rect 32204 62096 32220 62160
rect 32284 62156 37740 62160
rect 32284 62100 34385 62156
rect 34441 62100 37275 62156
rect 37331 62100 37740 62156
rect 32284 62096 37740 62100
rect 37804 62096 37820 62160
rect 37884 62096 37900 62160
rect 37964 62096 37980 62160
rect 38044 62096 38060 62160
rect 38124 62096 38140 62160
rect 38204 62096 38220 62160
rect 38284 62156 43740 62160
rect 38284 62100 40165 62156
rect 40221 62100 43055 62156
rect 43111 62100 43740 62156
rect 38284 62096 43740 62100
rect 43804 62096 43820 62160
rect 43884 62096 43900 62160
rect 43964 62096 43980 62160
rect 44044 62096 44060 62160
rect 44124 62096 44140 62160
rect 44204 62096 44220 62160
rect 44284 62156 49740 62160
rect 49804 62156 49820 62160
rect 49884 62156 49900 62160
rect 44284 62100 45945 62156
rect 46001 62100 48892 62156
rect 48948 62100 49740 62156
rect 49810 62100 49820 62156
rect 49890 62100 49900 62156
rect 44284 62096 49740 62100
rect 49804 62096 49820 62100
rect 49884 62096 49900 62100
rect 49964 62096 49980 62160
rect 50044 62096 50060 62160
rect 50124 62096 50140 62160
rect 50204 62096 50220 62160
rect 50284 62156 55740 62160
rect 50284 62100 53048 62156
rect 53104 62100 53206 62156
rect 53262 62100 53562 62156
rect 53618 62100 54880 62156
rect 54936 62100 55473 62156
rect 55529 62100 55740 62156
rect 50284 62096 55740 62100
rect 55804 62096 55820 62160
rect 55884 62096 55900 62160
rect 55964 62096 55980 62160
rect 56044 62096 56060 62160
rect 56124 62096 56140 62160
rect 56204 62096 56220 62160
rect 56284 62156 61740 62160
rect 56284 62100 56619 62156
rect 56675 62100 58055 62156
rect 58111 62100 58135 62156
rect 58191 62100 59298 62156
rect 59354 62100 59456 62156
rect 59512 62100 59764 62156
rect 59820 62100 59910 62156
rect 59966 62100 60046 62156
rect 60102 62100 60126 62156
rect 60182 62100 61740 62156
rect 56284 62096 61740 62100
rect 61804 62096 61820 62160
rect 61884 62096 61900 62160
rect 61964 62096 61980 62160
rect 62044 62096 62060 62160
rect 62124 62096 62140 62160
rect 62204 62096 62220 62160
rect 62284 62156 67740 62160
rect 62284 62100 62418 62156
rect 62474 62100 62498 62156
rect 62554 62100 67740 62156
rect 62284 62096 67740 62100
rect 67804 62096 67820 62160
rect 67884 62096 67900 62160
rect 67964 62096 67980 62160
rect 68044 62096 68060 62160
rect 68124 62096 68140 62160
rect 68204 62096 68220 62160
rect 68284 62156 73740 62160
rect 68284 62100 71864 62156
rect 71920 62100 71944 62156
rect 72000 62100 72024 62156
rect 72080 62100 72104 62156
rect 72160 62100 73740 62156
rect 68284 62096 73740 62100
rect 73804 62096 73820 62160
rect 73884 62096 73900 62160
rect 73964 62096 73980 62160
rect 74044 62096 74060 62160
rect 74124 62096 74140 62160
rect 74204 62096 74220 62160
rect 74284 62096 75028 62160
rect 964 62080 75028 62096
rect 964 62016 1740 62080
rect 1804 62016 1820 62080
rect 1884 62016 1900 62080
rect 1964 62016 1980 62080
rect 2044 62016 2060 62080
rect 2124 62016 2140 62080
rect 2204 62016 2220 62080
rect 2284 62076 7740 62080
rect 2332 62020 2356 62076
rect 2412 62020 5485 62076
rect 5541 62020 7740 62076
rect 2284 62016 7740 62020
rect 7804 62016 7820 62080
rect 7884 62016 7900 62080
rect 7964 62016 7980 62080
rect 8044 62016 8060 62080
rect 8124 62016 8140 62080
rect 8204 62016 8220 62080
rect 8284 62076 13740 62080
rect 8284 62020 8375 62076
rect 8431 62020 11265 62076
rect 11321 62020 13740 62076
rect 8284 62016 13740 62020
rect 13804 62016 13820 62080
rect 13884 62016 13900 62080
rect 13964 62016 13980 62080
rect 14044 62016 14060 62080
rect 14124 62016 14140 62080
rect 14204 62076 14220 62080
rect 14211 62020 14220 62076
rect 14204 62016 14220 62020
rect 14284 62076 19740 62080
rect 14284 62020 17045 62076
rect 17101 62020 19740 62076
rect 14284 62016 19740 62020
rect 19804 62016 19820 62080
rect 19884 62016 19900 62080
rect 19964 62076 19980 62080
rect 19964 62016 19980 62020
rect 20044 62016 20060 62080
rect 20124 62016 20140 62080
rect 20204 62016 20220 62080
rect 20284 62076 25740 62080
rect 20284 62020 22825 62076
rect 22881 62020 25715 62076
rect 20284 62016 25740 62020
rect 25804 62016 25820 62080
rect 25884 62016 25900 62080
rect 25964 62016 25980 62080
rect 26044 62016 26060 62080
rect 26124 62016 26140 62080
rect 26204 62016 26220 62080
rect 26284 62076 31740 62080
rect 26284 62020 28605 62076
rect 28661 62020 31495 62076
rect 31551 62020 31740 62076
rect 26284 62016 31740 62020
rect 31804 62016 31820 62080
rect 31884 62016 31900 62080
rect 31964 62016 31980 62080
rect 32044 62016 32060 62080
rect 32124 62016 32140 62080
rect 32204 62016 32220 62080
rect 32284 62076 37740 62080
rect 32284 62020 34385 62076
rect 34441 62020 37275 62076
rect 37331 62020 37740 62076
rect 32284 62016 37740 62020
rect 37804 62016 37820 62080
rect 37884 62016 37900 62080
rect 37964 62016 37980 62080
rect 38044 62016 38060 62080
rect 38124 62016 38140 62080
rect 38204 62016 38220 62080
rect 38284 62076 43740 62080
rect 38284 62020 40165 62076
rect 40221 62020 43055 62076
rect 43111 62020 43740 62076
rect 38284 62016 43740 62020
rect 43804 62016 43820 62080
rect 43884 62016 43900 62080
rect 43964 62016 43980 62080
rect 44044 62016 44060 62080
rect 44124 62016 44140 62080
rect 44204 62016 44220 62080
rect 44284 62076 49740 62080
rect 49804 62076 49820 62080
rect 49884 62076 49900 62080
rect 44284 62020 45945 62076
rect 46001 62020 48892 62076
rect 48948 62020 49740 62076
rect 49810 62020 49820 62076
rect 49890 62020 49900 62076
rect 44284 62016 49740 62020
rect 49804 62016 49820 62020
rect 49884 62016 49900 62020
rect 49964 62016 49980 62080
rect 50044 62016 50060 62080
rect 50124 62016 50140 62080
rect 50204 62016 50220 62080
rect 50284 62076 55740 62080
rect 50284 62020 53048 62076
rect 53104 62020 53206 62076
rect 53262 62020 53562 62076
rect 53618 62020 54880 62076
rect 54936 62020 55473 62076
rect 55529 62020 55740 62076
rect 50284 62016 55740 62020
rect 55804 62016 55820 62080
rect 55884 62016 55900 62080
rect 55964 62016 55980 62080
rect 56044 62016 56060 62080
rect 56124 62016 56140 62080
rect 56204 62016 56220 62080
rect 56284 62076 61740 62080
rect 56284 62020 56619 62076
rect 56675 62020 58055 62076
rect 58111 62020 58135 62076
rect 58191 62020 59298 62076
rect 59354 62020 59456 62076
rect 59512 62020 59764 62076
rect 59820 62020 59910 62076
rect 59966 62020 60046 62076
rect 60102 62020 60126 62076
rect 60182 62020 61740 62076
rect 56284 62016 61740 62020
rect 61804 62016 61820 62080
rect 61884 62016 61900 62080
rect 61964 62016 61980 62080
rect 62044 62016 62060 62080
rect 62124 62016 62140 62080
rect 62204 62016 62220 62080
rect 62284 62076 67740 62080
rect 62284 62020 62418 62076
rect 62474 62020 62498 62076
rect 62554 62020 67740 62076
rect 62284 62016 67740 62020
rect 67804 62016 67820 62080
rect 67884 62016 67900 62080
rect 67964 62016 67980 62080
rect 68044 62016 68060 62080
rect 68124 62016 68140 62080
rect 68204 62016 68220 62080
rect 68284 62076 73740 62080
rect 68284 62020 71864 62076
rect 71920 62020 71944 62076
rect 72000 62020 72024 62076
rect 72080 62020 72104 62076
rect 72160 62020 73740 62076
rect 68284 62016 73740 62020
rect 73804 62016 73820 62080
rect 73884 62016 73900 62080
rect 73964 62016 73980 62080
rect 74044 62016 74060 62080
rect 74124 62016 74140 62080
rect 74204 62016 74220 62080
rect 74284 62016 75028 62080
rect 964 62000 75028 62016
rect 964 61936 1740 62000
rect 1804 61936 1820 62000
rect 1884 61936 1900 62000
rect 1964 61936 1980 62000
rect 2044 61936 2060 62000
rect 2124 61936 2140 62000
rect 2204 61936 2220 62000
rect 2284 61996 7740 62000
rect 2332 61940 2356 61996
rect 2412 61940 5485 61996
rect 5541 61940 7740 61996
rect 2284 61936 7740 61940
rect 7804 61936 7820 62000
rect 7884 61936 7900 62000
rect 7964 61936 7980 62000
rect 8044 61936 8060 62000
rect 8124 61936 8140 62000
rect 8204 61936 8220 62000
rect 8284 61996 13740 62000
rect 8284 61940 8375 61996
rect 8431 61940 11265 61996
rect 11321 61940 13740 61996
rect 8284 61936 13740 61940
rect 13804 61936 13820 62000
rect 13884 61936 13900 62000
rect 13964 61936 13980 62000
rect 14044 61936 14060 62000
rect 14124 61936 14140 62000
rect 14204 61996 14220 62000
rect 14211 61940 14220 61996
rect 14204 61936 14220 61940
rect 14284 61996 19740 62000
rect 14284 61940 17045 61996
rect 17101 61940 19740 61996
rect 14284 61936 19740 61940
rect 19804 61936 19820 62000
rect 19884 61936 19900 62000
rect 19964 61996 19980 62000
rect 19964 61936 19980 61940
rect 20044 61936 20060 62000
rect 20124 61936 20140 62000
rect 20204 61936 20220 62000
rect 20284 61996 25740 62000
rect 20284 61940 22825 61996
rect 22881 61940 25715 61996
rect 20284 61936 25740 61940
rect 25804 61936 25820 62000
rect 25884 61936 25900 62000
rect 25964 61936 25980 62000
rect 26044 61936 26060 62000
rect 26124 61936 26140 62000
rect 26204 61936 26220 62000
rect 26284 61996 31740 62000
rect 26284 61940 28605 61996
rect 28661 61940 31495 61996
rect 31551 61940 31740 61996
rect 26284 61936 31740 61940
rect 31804 61936 31820 62000
rect 31884 61936 31900 62000
rect 31964 61936 31980 62000
rect 32044 61936 32060 62000
rect 32124 61936 32140 62000
rect 32204 61936 32220 62000
rect 32284 61996 37740 62000
rect 32284 61940 34385 61996
rect 34441 61940 37275 61996
rect 37331 61940 37740 61996
rect 32284 61936 37740 61940
rect 37804 61936 37820 62000
rect 37884 61936 37900 62000
rect 37964 61936 37980 62000
rect 38044 61936 38060 62000
rect 38124 61936 38140 62000
rect 38204 61936 38220 62000
rect 38284 61996 43740 62000
rect 38284 61940 40165 61996
rect 40221 61940 43055 61996
rect 43111 61940 43740 61996
rect 38284 61936 43740 61940
rect 43804 61936 43820 62000
rect 43884 61936 43900 62000
rect 43964 61936 43980 62000
rect 44044 61936 44060 62000
rect 44124 61936 44140 62000
rect 44204 61936 44220 62000
rect 44284 61996 49740 62000
rect 49804 61996 49820 62000
rect 49884 61996 49900 62000
rect 44284 61940 45945 61996
rect 46001 61940 48892 61996
rect 48948 61940 49740 61996
rect 49810 61940 49820 61996
rect 49890 61940 49900 61996
rect 44284 61936 49740 61940
rect 49804 61936 49820 61940
rect 49884 61936 49900 61940
rect 49964 61936 49980 62000
rect 50044 61936 50060 62000
rect 50124 61936 50140 62000
rect 50204 61936 50220 62000
rect 50284 61996 55740 62000
rect 50284 61940 53048 61996
rect 53104 61940 53206 61996
rect 53262 61940 53562 61996
rect 53618 61940 54880 61996
rect 54936 61940 55473 61996
rect 55529 61940 55740 61996
rect 50284 61936 55740 61940
rect 55804 61936 55820 62000
rect 55884 61936 55900 62000
rect 55964 61936 55980 62000
rect 56044 61936 56060 62000
rect 56124 61936 56140 62000
rect 56204 61936 56220 62000
rect 56284 61996 61740 62000
rect 56284 61940 56619 61996
rect 56675 61940 58055 61996
rect 58111 61940 58135 61996
rect 58191 61940 59298 61996
rect 59354 61940 59456 61996
rect 59512 61940 59764 61996
rect 59820 61940 59910 61996
rect 59966 61940 60046 61996
rect 60102 61940 60126 61996
rect 60182 61940 61740 61996
rect 56284 61936 61740 61940
rect 61804 61936 61820 62000
rect 61884 61936 61900 62000
rect 61964 61936 61980 62000
rect 62044 61936 62060 62000
rect 62124 61936 62140 62000
rect 62204 61936 62220 62000
rect 62284 61996 67740 62000
rect 62284 61940 62418 61996
rect 62474 61940 62498 61996
rect 62554 61940 67740 61996
rect 62284 61936 67740 61940
rect 67804 61936 67820 62000
rect 67884 61936 67900 62000
rect 67964 61936 67980 62000
rect 68044 61936 68060 62000
rect 68124 61936 68140 62000
rect 68204 61936 68220 62000
rect 68284 61996 73740 62000
rect 68284 61940 71864 61996
rect 71920 61940 71944 61996
rect 72000 61940 72024 61996
rect 72080 61940 72104 61996
rect 72160 61940 73740 61996
rect 68284 61936 73740 61940
rect 73804 61936 73820 62000
rect 73884 61936 73900 62000
rect 73964 61936 73980 62000
rect 74044 61936 74060 62000
rect 74124 61936 74140 62000
rect 74204 61936 74220 62000
rect 74284 61936 75028 62000
rect 964 61912 75028 61936
rect 63493 61026 63559 61029
rect 63902 61026 63908 61028
rect 63493 61024 63908 61026
rect 63493 60968 63498 61024
rect 63554 60968 63908 61024
rect 63493 60966 63908 60968
rect 63493 60963 63559 60966
rect 63902 60964 63908 60966
rect 63972 60964 63978 61028
rect 63493 58714 63559 58717
rect 64086 58714 64092 58716
rect 63493 58712 64092 58714
rect 63493 58656 63498 58712
rect 63554 58656 64092 58712
rect 63493 58654 64092 58656
rect 63493 58651 63559 58654
rect 64086 58652 64092 58654
rect 64156 58652 64162 58716
rect 63493 56674 63559 56677
rect 64270 56674 64276 56676
rect 63493 56672 64276 56674
rect 63493 56616 63498 56672
rect 63554 56616 64276 56672
rect 63493 56614 64276 56616
rect 63493 56611 63559 56614
rect 64270 56612 64276 56614
rect 64340 56612 64346 56676
rect 63493 54770 63559 54773
rect 69054 54770 69060 54772
rect 63493 54768 69060 54770
rect 63493 54712 63498 54768
rect 63554 54712 69060 54768
rect 63493 54710 69060 54712
rect 63493 54707 63559 54710
rect 69054 54708 69060 54710
rect 69124 54708 69130 54772
rect 964 54592 75028 54616
rect 964 54588 4740 54592
rect 964 54532 2136 54588
rect 2192 54532 4740 54588
rect 964 54528 4740 54532
rect 4804 54528 4820 54592
rect 4884 54528 4900 54592
rect 4964 54528 4980 54592
rect 5044 54528 5060 54592
rect 5124 54528 5140 54592
rect 5204 54528 5220 54592
rect 5284 54588 10740 54592
rect 5284 54532 5632 54588
rect 5688 54532 8522 54588
rect 8578 54532 10740 54588
rect 5284 54528 10740 54532
rect 10804 54528 10820 54592
rect 10884 54528 10900 54592
rect 10964 54528 10980 54592
rect 11044 54528 11060 54592
rect 11124 54528 11140 54592
rect 11204 54528 11220 54592
rect 11284 54588 16740 54592
rect 11284 54532 11412 54588
rect 11468 54532 14302 54588
rect 14358 54532 16740 54588
rect 11284 54528 16740 54532
rect 16804 54528 16820 54592
rect 16884 54528 16900 54592
rect 16964 54528 16980 54592
rect 17044 54528 17060 54592
rect 17124 54528 17140 54592
rect 17204 54588 17220 54592
rect 17284 54588 22740 54592
rect 17284 54532 20082 54588
rect 20138 54532 22740 54588
rect 17204 54528 17220 54532
rect 17284 54528 22740 54532
rect 22804 54528 22820 54592
rect 22884 54528 22900 54592
rect 22964 54588 22980 54592
rect 22964 54532 22972 54588
rect 22964 54528 22980 54532
rect 23044 54528 23060 54592
rect 23124 54528 23140 54592
rect 23204 54528 23220 54592
rect 23284 54588 28740 54592
rect 28804 54588 28820 54592
rect 23284 54532 25862 54588
rect 25918 54532 28740 54588
rect 28808 54532 28820 54588
rect 23284 54528 28740 54532
rect 28804 54528 28820 54532
rect 28884 54528 28900 54592
rect 28964 54528 28980 54592
rect 29044 54528 29060 54592
rect 29124 54528 29140 54592
rect 29204 54528 29220 54592
rect 29284 54588 34740 54592
rect 29284 54532 31642 54588
rect 31698 54532 34532 54588
rect 34588 54532 34740 54588
rect 29284 54528 34740 54532
rect 34804 54528 34820 54592
rect 34884 54528 34900 54592
rect 34964 54528 34980 54592
rect 35044 54528 35060 54592
rect 35124 54528 35140 54592
rect 35204 54528 35220 54592
rect 35284 54588 40740 54592
rect 35284 54532 37422 54588
rect 37478 54532 40312 54588
rect 40368 54532 40740 54588
rect 35284 54528 40740 54532
rect 40804 54528 40820 54592
rect 40884 54528 40900 54592
rect 40964 54528 40980 54592
rect 41044 54528 41060 54592
rect 41124 54528 41140 54592
rect 41204 54528 41220 54592
rect 41284 54588 46740 54592
rect 41284 54532 43202 54588
rect 43258 54532 46092 54588
rect 46148 54532 46740 54588
rect 41284 54528 46740 54532
rect 46804 54528 46820 54592
rect 46884 54528 46900 54592
rect 46964 54528 46980 54592
rect 47044 54528 47060 54592
rect 47124 54528 47140 54592
rect 47204 54528 47220 54592
rect 47284 54588 52740 54592
rect 47284 54532 49100 54588
rect 49156 54532 52329 54588
rect 52385 54532 52740 54588
rect 47284 54528 52740 54532
rect 52804 54528 52820 54592
rect 52884 54528 52900 54592
rect 52964 54528 52980 54592
rect 53044 54528 53060 54592
rect 53124 54528 53140 54592
rect 53204 54528 53220 54592
rect 53284 54588 58740 54592
rect 53284 54532 53730 54588
rect 53786 54532 53898 54588
rect 53954 54532 54642 54588
rect 54698 54532 55032 54588
rect 55088 54532 55748 54588
rect 55804 54532 56326 54588
rect 56382 54532 56771 54588
rect 56827 54532 57075 54588
rect 57131 54532 57917 54588
rect 57973 54532 58557 54588
rect 58613 54532 58740 54588
rect 53284 54528 58740 54532
rect 58804 54528 58820 54592
rect 58884 54528 58900 54592
rect 58964 54528 58980 54592
rect 59044 54528 59060 54592
rect 59124 54528 59140 54592
rect 59204 54528 59220 54592
rect 59284 54588 64740 54592
rect 59284 54532 60418 54588
rect 60474 54532 60576 54588
rect 60632 54532 62620 54588
rect 62676 54532 62700 54588
rect 62756 54532 64740 54588
rect 59284 54528 64740 54532
rect 64804 54528 64820 54592
rect 64884 54528 64900 54592
rect 64964 54528 64980 54592
rect 65044 54528 65060 54592
rect 65124 54528 65140 54592
rect 65204 54528 65220 54592
rect 65284 54528 70740 54592
rect 70804 54528 70820 54592
rect 70884 54528 70900 54592
rect 70964 54528 70980 54592
rect 71044 54528 71060 54592
rect 71124 54528 71140 54592
rect 71204 54528 71220 54592
rect 71284 54588 75028 54592
rect 71284 54532 74216 54588
rect 74272 54532 74296 54588
rect 74352 54532 74376 54588
rect 74432 54532 74456 54588
rect 74512 54532 75028 54588
rect 71284 54528 75028 54532
rect 964 54512 75028 54528
rect 964 54508 4740 54512
rect 964 54452 2136 54508
rect 2192 54452 4740 54508
rect 964 54448 4740 54452
rect 4804 54448 4820 54512
rect 4884 54448 4900 54512
rect 4964 54448 4980 54512
rect 5044 54448 5060 54512
rect 5124 54448 5140 54512
rect 5204 54448 5220 54512
rect 5284 54508 10740 54512
rect 5284 54452 5632 54508
rect 5688 54452 8522 54508
rect 8578 54452 10740 54508
rect 5284 54448 10740 54452
rect 10804 54448 10820 54512
rect 10884 54448 10900 54512
rect 10964 54448 10980 54512
rect 11044 54448 11060 54512
rect 11124 54448 11140 54512
rect 11204 54448 11220 54512
rect 11284 54508 16740 54512
rect 11284 54452 11412 54508
rect 11468 54452 14302 54508
rect 14358 54452 16740 54508
rect 11284 54448 16740 54452
rect 16804 54448 16820 54512
rect 16884 54448 16900 54512
rect 16964 54448 16980 54512
rect 17044 54448 17060 54512
rect 17124 54448 17140 54512
rect 17204 54508 17220 54512
rect 17284 54508 22740 54512
rect 17284 54452 20082 54508
rect 20138 54452 22740 54508
rect 17204 54448 17220 54452
rect 17284 54448 22740 54452
rect 22804 54448 22820 54512
rect 22884 54448 22900 54512
rect 22964 54508 22980 54512
rect 22964 54452 22972 54508
rect 22964 54448 22980 54452
rect 23044 54448 23060 54512
rect 23124 54448 23140 54512
rect 23204 54448 23220 54512
rect 23284 54508 28740 54512
rect 28804 54508 28820 54512
rect 23284 54452 25862 54508
rect 25918 54452 28740 54508
rect 28808 54452 28820 54508
rect 23284 54448 28740 54452
rect 28804 54448 28820 54452
rect 28884 54448 28900 54512
rect 28964 54448 28980 54512
rect 29044 54448 29060 54512
rect 29124 54448 29140 54512
rect 29204 54448 29220 54512
rect 29284 54508 34740 54512
rect 29284 54452 31642 54508
rect 31698 54452 34532 54508
rect 34588 54452 34740 54508
rect 29284 54448 34740 54452
rect 34804 54448 34820 54512
rect 34884 54448 34900 54512
rect 34964 54448 34980 54512
rect 35044 54448 35060 54512
rect 35124 54448 35140 54512
rect 35204 54448 35220 54512
rect 35284 54508 40740 54512
rect 35284 54452 37422 54508
rect 37478 54452 40312 54508
rect 40368 54452 40740 54508
rect 35284 54448 40740 54452
rect 40804 54448 40820 54512
rect 40884 54448 40900 54512
rect 40964 54448 40980 54512
rect 41044 54448 41060 54512
rect 41124 54448 41140 54512
rect 41204 54448 41220 54512
rect 41284 54508 46740 54512
rect 41284 54452 43202 54508
rect 43258 54452 46092 54508
rect 46148 54452 46740 54508
rect 41284 54448 46740 54452
rect 46804 54448 46820 54512
rect 46884 54448 46900 54512
rect 46964 54448 46980 54512
rect 47044 54448 47060 54512
rect 47124 54448 47140 54512
rect 47204 54448 47220 54512
rect 47284 54508 52740 54512
rect 47284 54452 49100 54508
rect 49156 54452 52329 54508
rect 52385 54452 52740 54508
rect 47284 54448 52740 54452
rect 52804 54448 52820 54512
rect 52884 54448 52900 54512
rect 52964 54448 52980 54512
rect 53044 54448 53060 54512
rect 53124 54448 53140 54512
rect 53204 54448 53220 54512
rect 53284 54508 58740 54512
rect 53284 54452 53730 54508
rect 53786 54452 53898 54508
rect 53954 54452 54642 54508
rect 54698 54452 55032 54508
rect 55088 54452 55748 54508
rect 55804 54452 56326 54508
rect 56382 54452 56771 54508
rect 56827 54452 57075 54508
rect 57131 54452 57917 54508
rect 57973 54452 58557 54508
rect 58613 54452 58740 54508
rect 53284 54448 58740 54452
rect 58804 54448 58820 54512
rect 58884 54448 58900 54512
rect 58964 54448 58980 54512
rect 59044 54448 59060 54512
rect 59124 54448 59140 54512
rect 59204 54448 59220 54512
rect 59284 54508 64740 54512
rect 59284 54452 60418 54508
rect 60474 54452 60576 54508
rect 60632 54452 62620 54508
rect 62676 54452 62700 54508
rect 62756 54452 64740 54508
rect 59284 54448 64740 54452
rect 64804 54448 64820 54512
rect 64884 54448 64900 54512
rect 64964 54448 64980 54512
rect 65044 54448 65060 54512
rect 65124 54448 65140 54512
rect 65204 54448 65220 54512
rect 65284 54448 70740 54512
rect 70804 54448 70820 54512
rect 70884 54448 70900 54512
rect 70964 54448 70980 54512
rect 71044 54448 71060 54512
rect 71124 54448 71140 54512
rect 71204 54448 71220 54512
rect 71284 54508 75028 54512
rect 71284 54452 74216 54508
rect 74272 54452 74296 54508
rect 74352 54452 74376 54508
rect 74432 54452 74456 54508
rect 74512 54452 75028 54508
rect 71284 54448 75028 54452
rect 964 54432 75028 54448
rect 964 54428 4740 54432
rect 964 54372 2136 54428
rect 2192 54372 4740 54428
rect 964 54368 4740 54372
rect 4804 54368 4820 54432
rect 4884 54368 4900 54432
rect 4964 54368 4980 54432
rect 5044 54368 5060 54432
rect 5124 54368 5140 54432
rect 5204 54368 5220 54432
rect 5284 54428 10740 54432
rect 5284 54372 5632 54428
rect 5688 54372 8522 54428
rect 8578 54372 10740 54428
rect 5284 54368 10740 54372
rect 10804 54368 10820 54432
rect 10884 54368 10900 54432
rect 10964 54368 10980 54432
rect 11044 54368 11060 54432
rect 11124 54368 11140 54432
rect 11204 54368 11220 54432
rect 11284 54428 16740 54432
rect 11284 54372 11412 54428
rect 11468 54372 14302 54428
rect 14358 54372 16740 54428
rect 11284 54368 16740 54372
rect 16804 54368 16820 54432
rect 16884 54368 16900 54432
rect 16964 54368 16980 54432
rect 17044 54368 17060 54432
rect 17124 54368 17140 54432
rect 17204 54428 17220 54432
rect 17284 54428 22740 54432
rect 17284 54372 20082 54428
rect 20138 54372 22740 54428
rect 17204 54368 17220 54372
rect 17284 54368 22740 54372
rect 22804 54368 22820 54432
rect 22884 54368 22900 54432
rect 22964 54428 22980 54432
rect 22964 54372 22972 54428
rect 22964 54368 22980 54372
rect 23044 54368 23060 54432
rect 23124 54368 23140 54432
rect 23204 54368 23220 54432
rect 23284 54428 28740 54432
rect 28804 54428 28820 54432
rect 23284 54372 25862 54428
rect 25918 54372 28740 54428
rect 28808 54372 28820 54428
rect 23284 54368 28740 54372
rect 28804 54368 28820 54372
rect 28884 54368 28900 54432
rect 28964 54368 28980 54432
rect 29044 54368 29060 54432
rect 29124 54368 29140 54432
rect 29204 54368 29220 54432
rect 29284 54428 34740 54432
rect 29284 54372 31642 54428
rect 31698 54372 34532 54428
rect 34588 54372 34740 54428
rect 29284 54368 34740 54372
rect 34804 54368 34820 54432
rect 34884 54368 34900 54432
rect 34964 54368 34980 54432
rect 35044 54368 35060 54432
rect 35124 54368 35140 54432
rect 35204 54368 35220 54432
rect 35284 54428 40740 54432
rect 35284 54372 37422 54428
rect 37478 54372 40312 54428
rect 40368 54372 40740 54428
rect 35284 54368 40740 54372
rect 40804 54368 40820 54432
rect 40884 54368 40900 54432
rect 40964 54368 40980 54432
rect 41044 54368 41060 54432
rect 41124 54368 41140 54432
rect 41204 54368 41220 54432
rect 41284 54428 46740 54432
rect 41284 54372 43202 54428
rect 43258 54372 46092 54428
rect 46148 54372 46740 54428
rect 41284 54368 46740 54372
rect 46804 54368 46820 54432
rect 46884 54368 46900 54432
rect 46964 54368 46980 54432
rect 47044 54368 47060 54432
rect 47124 54368 47140 54432
rect 47204 54368 47220 54432
rect 47284 54428 52740 54432
rect 47284 54372 49100 54428
rect 49156 54372 52329 54428
rect 52385 54372 52740 54428
rect 47284 54368 52740 54372
rect 52804 54368 52820 54432
rect 52884 54368 52900 54432
rect 52964 54368 52980 54432
rect 53044 54368 53060 54432
rect 53124 54368 53140 54432
rect 53204 54368 53220 54432
rect 53284 54428 58740 54432
rect 53284 54372 53730 54428
rect 53786 54372 53898 54428
rect 53954 54372 54642 54428
rect 54698 54372 55032 54428
rect 55088 54372 55748 54428
rect 55804 54372 56326 54428
rect 56382 54372 56771 54428
rect 56827 54372 57075 54428
rect 57131 54372 57917 54428
rect 57973 54372 58557 54428
rect 58613 54372 58740 54428
rect 53284 54368 58740 54372
rect 58804 54368 58820 54432
rect 58884 54368 58900 54432
rect 58964 54368 58980 54432
rect 59044 54368 59060 54432
rect 59124 54368 59140 54432
rect 59204 54368 59220 54432
rect 59284 54428 64740 54432
rect 59284 54372 60418 54428
rect 60474 54372 60576 54428
rect 60632 54372 62620 54428
rect 62676 54372 62700 54428
rect 62756 54372 64740 54428
rect 59284 54368 64740 54372
rect 64804 54368 64820 54432
rect 64884 54368 64900 54432
rect 64964 54368 64980 54432
rect 65044 54368 65060 54432
rect 65124 54368 65140 54432
rect 65204 54368 65220 54432
rect 65284 54368 70740 54432
rect 70804 54368 70820 54432
rect 70884 54368 70900 54432
rect 70964 54368 70980 54432
rect 71044 54368 71060 54432
rect 71124 54368 71140 54432
rect 71204 54368 71220 54432
rect 71284 54428 75028 54432
rect 71284 54372 74216 54428
rect 74272 54372 74296 54428
rect 74352 54372 74376 54428
rect 74432 54372 74456 54428
rect 74512 54372 75028 54428
rect 71284 54368 75028 54372
rect 964 54352 75028 54368
rect 964 54348 4740 54352
rect 964 54292 2136 54348
rect 2192 54292 4740 54348
rect 964 54288 4740 54292
rect 4804 54288 4820 54352
rect 4884 54288 4900 54352
rect 4964 54288 4980 54352
rect 5044 54288 5060 54352
rect 5124 54288 5140 54352
rect 5204 54288 5220 54352
rect 5284 54348 10740 54352
rect 5284 54292 5632 54348
rect 5688 54292 8522 54348
rect 8578 54292 10740 54348
rect 5284 54288 10740 54292
rect 10804 54288 10820 54352
rect 10884 54288 10900 54352
rect 10964 54288 10980 54352
rect 11044 54288 11060 54352
rect 11124 54288 11140 54352
rect 11204 54288 11220 54352
rect 11284 54348 16740 54352
rect 11284 54292 11412 54348
rect 11468 54292 14302 54348
rect 14358 54292 16740 54348
rect 11284 54288 16740 54292
rect 16804 54288 16820 54352
rect 16884 54288 16900 54352
rect 16964 54288 16980 54352
rect 17044 54288 17060 54352
rect 17124 54288 17140 54352
rect 17204 54348 17220 54352
rect 17284 54348 22740 54352
rect 17284 54292 20082 54348
rect 20138 54292 22740 54348
rect 17204 54288 17220 54292
rect 17284 54288 22740 54292
rect 22804 54288 22820 54352
rect 22884 54288 22900 54352
rect 22964 54348 22980 54352
rect 22964 54292 22972 54348
rect 22964 54288 22980 54292
rect 23044 54288 23060 54352
rect 23124 54288 23140 54352
rect 23204 54288 23220 54352
rect 23284 54348 28740 54352
rect 28804 54348 28820 54352
rect 23284 54292 25862 54348
rect 25918 54292 28740 54348
rect 28808 54292 28820 54348
rect 23284 54288 28740 54292
rect 28804 54288 28820 54292
rect 28884 54288 28900 54352
rect 28964 54288 28980 54352
rect 29044 54288 29060 54352
rect 29124 54288 29140 54352
rect 29204 54288 29220 54352
rect 29284 54348 34740 54352
rect 29284 54292 31642 54348
rect 31698 54292 34532 54348
rect 34588 54292 34740 54348
rect 29284 54288 34740 54292
rect 34804 54288 34820 54352
rect 34884 54288 34900 54352
rect 34964 54288 34980 54352
rect 35044 54288 35060 54352
rect 35124 54288 35140 54352
rect 35204 54288 35220 54352
rect 35284 54348 40740 54352
rect 35284 54292 37422 54348
rect 37478 54292 40312 54348
rect 40368 54292 40740 54348
rect 35284 54288 40740 54292
rect 40804 54288 40820 54352
rect 40884 54288 40900 54352
rect 40964 54288 40980 54352
rect 41044 54288 41060 54352
rect 41124 54288 41140 54352
rect 41204 54288 41220 54352
rect 41284 54348 46740 54352
rect 41284 54292 43202 54348
rect 43258 54292 46092 54348
rect 46148 54292 46740 54348
rect 41284 54288 46740 54292
rect 46804 54288 46820 54352
rect 46884 54288 46900 54352
rect 46964 54288 46980 54352
rect 47044 54288 47060 54352
rect 47124 54288 47140 54352
rect 47204 54288 47220 54352
rect 47284 54348 52740 54352
rect 47284 54292 49100 54348
rect 49156 54292 52329 54348
rect 52385 54292 52740 54348
rect 47284 54288 52740 54292
rect 52804 54288 52820 54352
rect 52884 54288 52900 54352
rect 52964 54288 52980 54352
rect 53044 54288 53060 54352
rect 53124 54288 53140 54352
rect 53204 54288 53220 54352
rect 53284 54348 58740 54352
rect 53284 54292 53730 54348
rect 53786 54292 53898 54348
rect 53954 54292 54642 54348
rect 54698 54292 55032 54348
rect 55088 54292 55748 54348
rect 55804 54292 56326 54348
rect 56382 54292 56771 54348
rect 56827 54292 57075 54348
rect 57131 54292 57917 54348
rect 57973 54292 58557 54348
rect 58613 54292 58740 54348
rect 53284 54288 58740 54292
rect 58804 54288 58820 54352
rect 58884 54288 58900 54352
rect 58964 54288 58980 54352
rect 59044 54288 59060 54352
rect 59124 54288 59140 54352
rect 59204 54288 59220 54352
rect 59284 54348 64740 54352
rect 59284 54292 60418 54348
rect 60474 54292 60576 54348
rect 60632 54292 62620 54348
rect 62676 54292 62700 54348
rect 62756 54292 64740 54348
rect 59284 54288 64740 54292
rect 64804 54288 64820 54352
rect 64884 54288 64900 54352
rect 64964 54288 64980 54352
rect 65044 54288 65060 54352
rect 65124 54288 65140 54352
rect 65204 54288 65220 54352
rect 65284 54288 70740 54352
rect 70804 54288 70820 54352
rect 70884 54288 70900 54352
rect 70964 54288 70980 54352
rect 71044 54288 71060 54352
rect 71124 54288 71140 54352
rect 71204 54288 71220 54352
rect 71284 54348 75028 54352
rect 71284 54292 74216 54348
rect 74272 54292 74296 54348
rect 74352 54292 74376 54348
rect 74432 54292 74456 54348
rect 74512 54292 75028 54348
rect 71284 54288 75028 54292
rect 964 54264 75028 54288
rect 964 52240 75028 52264
rect 964 52176 1740 52240
rect 1804 52176 1820 52240
rect 1884 52176 1900 52240
rect 1964 52176 1980 52240
rect 2044 52176 2060 52240
rect 2124 52176 2140 52240
rect 2204 52176 2220 52240
rect 2284 52236 7740 52240
rect 2332 52180 2356 52236
rect 2412 52180 5485 52236
rect 5541 52180 7740 52236
rect 2284 52176 7740 52180
rect 7804 52176 7820 52240
rect 7884 52176 7900 52240
rect 7964 52176 7980 52240
rect 8044 52176 8060 52240
rect 8124 52176 8140 52240
rect 8204 52176 8220 52240
rect 8284 52236 13740 52240
rect 8284 52180 8375 52236
rect 8431 52180 11265 52236
rect 11321 52180 13740 52236
rect 8284 52176 13740 52180
rect 13804 52176 13820 52240
rect 13884 52176 13900 52240
rect 13964 52176 13980 52240
rect 14044 52176 14060 52240
rect 14124 52176 14140 52240
rect 14204 52236 14220 52240
rect 14211 52180 14220 52236
rect 14204 52176 14220 52180
rect 14284 52236 19740 52240
rect 14284 52180 17045 52236
rect 17101 52180 19740 52236
rect 14284 52176 19740 52180
rect 19804 52176 19820 52240
rect 19884 52176 19900 52240
rect 19964 52236 19980 52240
rect 19964 52176 19980 52180
rect 20044 52176 20060 52240
rect 20124 52176 20140 52240
rect 20204 52176 20220 52240
rect 20284 52236 25740 52240
rect 20284 52180 22825 52236
rect 22881 52180 25715 52236
rect 20284 52176 25740 52180
rect 25804 52176 25820 52240
rect 25884 52176 25900 52240
rect 25964 52176 25980 52240
rect 26044 52176 26060 52240
rect 26124 52176 26140 52240
rect 26204 52176 26220 52240
rect 26284 52236 31740 52240
rect 26284 52180 28605 52236
rect 28661 52180 31495 52236
rect 31551 52180 31740 52236
rect 26284 52176 31740 52180
rect 31804 52176 31820 52240
rect 31884 52176 31900 52240
rect 31964 52176 31980 52240
rect 32044 52176 32060 52240
rect 32124 52176 32140 52240
rect 32204 52176 32220 52240
rect 32284 52236 37740 52240
rect 32284 52180 34385 52236
rect 34441 52180 37275 52236
rect 37331 52180 37740 52236
rect 32284 52176 37740 52180
rect 37804 52176 37820 52240
rect 37884 52176 37900 52240
rect 37964 52176 37980 52240
rect 38044 52176 38060 52240
rect 38124 52176 38140 52240
rect 38204 52176 38220 52240
rect 38284 52236 43740 52240
rect 38284 52180 40165 52236
rect 40221 52180 43055 52236
rect 43111 52180 43740 52236
rect 38284 52176 43740 52180
rect 43804 52176 43820 52240
rect 43884 52176 43900 52240
rect 43964 52176 43980 52240
rect 44044 52176 44060 52240
rect 44124 52176 44140 52240
rect 44204 52176 44220 52240
rect 44284 52236 49740 52240
rect 49804 52236 49820 52240
rect 49884 52236 49900 52240
rect 44284 52180 45945 52236
rect 46001 52180 48892 52236
rect 48948 52180 49740 52236
rect 49810 52180 49820 52236
rect 49890 52180 49900 52236
rect 44284 52176 49740 52180
rect 49804 52176 49820 52180
rect 49884 52176 49900 52180
rect 49964 52176 49980 52240
rect 50044 52176 50060 52240
rect 50124 52176 50140 52240
rect 50204 52176 50220 52240
rect 50284 52236 55740 52240
rect 50284 52180 53048 52236
rect 53104 52180 53206 52236
rect 53262 52180 53562 52236
rect 53618 52180 54880 52236
rect 54936 52180 55473 52236
rect 55529 52180 55740 52236
rect 50284 52176 55740 52180
rect 55804 52176 55820 52240
rect 55884 52176 55900 52240
rect 55964 52176 55980 52240
rect 56044 52176 56060 52240
rect 56124 52176 56140 52240
rect 56204 52176 56220 52240
rect 56284 52236 61740 52240
rect 56284 52180 56619 52236
rect 56675 52180 58055 52236
rect 58111 52180 58135 52236
rect 58191 52180 59298 52236
rect 59354 52180 59456 52236
rect 59512 52180 59764 52236
rect 59820 52180 59910 52236
rect 59966 52180 60046 52236
rect 60102 52180 60126 52236
rect 60182 52180 61740 52236
rect 56284 52176 61740 52180
rect 61804 52176 61820 52240
rect 61884 52176 61900 52240
rect 61964 52176 61980 52240
rect 62044 52176 62060 52240
rect 62124 52176 62140 52240
rect 62204 52176 62220 52240
rect 62284 52236 67740 52240
rect 62284 52180 62418 52236
rect 62474 52180 62498 52236
rect 62554 52180 67740 52236
rect 62284 52176 67740 52180
rect 67804 52176 67820 52240
rect 67884 52176 67900 52240
rect 67964 52176 67980 52240
rect 68044 52176 68060 52240
rect 68124 52176 68140 52240
rect 68204 52176 68220 52240
rect 68284 52236 73740 52240
rect 68284 52180 71864 52236
rect 71920 52180 71944 52236
rect 72000 52180 72024 52236
rect 72080 52180 72104 52236
rect 72160 52180 73740 52236
rect 68284 52176 73740 52180
rect 73804 52176 73820 52240
rect 73884 52176 73900 52240
rect 73964 52176 73980 52240
rect 74044 52176 74060 52240
rect 74124 52176 74140 52240
rect 74204 52176 74220 52240
rect 74284 52176 75028 52240
rect 964 52160 75028 52176
rect 964 52096 1740 52160
rect 1804 52096 1820 52160
rect 1884 52096 1900 52160
rect 1964 52096 1980 52160
rect 2044 52096 2060 52160
rect 2124 52096 2140 52160
rect 2204 52096 2220 52160
rect 2284 52156 7740 52160
rect 2332 52100 2356 52156
rect 2412 52100 5485 52156
rect 5541 52100 7740 52156
rect 2284 52096 7740 52100
rect 7804 52096 7820 52160
rect 7884 52096 7900 52160
rect 7964 52096 7980 52160
rect 8044 52096 8060 52160
rect 8124 52096 8140 52160
rect 8204 52096 8220 52160
rect 8284 52156 13740 52160
rect 8284 52100 8375 52156
rect 8431 52100 11265 52156
rect 11321 52100 13740 52156
rect 8284 52096 13740 52100
rect 13804 52096 13820 52160
rect 13884 52096 13900 52160
rect 13964 52096 13980 52160
rect 14044 52096 14060 52160
rect 14124 52096 14140 52160
rect 14204 52156 14220 52160
rect 14211 52100 14220 52156
rect 14204 52096 14220 52100
rect 14284 52156 19740 52160
rect 14284 52100 17045 52156
rect 17101 52100 19740 52156
rect 14284 52096 19740 52100
rect 19804 52096 19820 52160
rect 19884 52096 19900 52160
rect 19964 52156 19980 52160
rect 19964 52096 19980 52100
rect 20044 52096 20060 52160
rect 20124 52096 20140 52160
rect 20204 52096 20220 52160
rect 20284 52156 25740 52160
rect 20284 52100 22825 52156
rect 22881 52100 25715 52156
rect 20284 52096 25740 52100
rect 25804 52096 25820 52160
rect 25884 52096 25900 52160
rect 25964 52096 25980 52160
rect 26044 52096 26060 52160
rect 26124 52096 26140 52160
rect 26204 52096 26220 52160
rect 26284 52156 31740 52160
rect 26284 52100 28605 52156
rect 28661 52100 31495 52156
rect 31551 52100 31740 52156
rect 26284 52096 31740 52100
rect 31804 52096 31820 52160
rect 31884 52096 31900 52160
rect 31964 52096 31980 52160
rect 32044 52096 32060 52160
rect 32124 52096 32140 52160
rect 32204 52096 32220 52160
rect 32284 52156 37740 52160
rect 32284 52100 34385 52156
rect 34441 52100 37275 52156
rect 37331 52100 37740 52156
rect 32284 52096 37740 52100
rect 37804 52096 37820 52160
rect 37884 52096 37900 52160
rect 37964 52096 37980 52160
rect 38044 52096 38060 52160
rect 38124 52096 38140 52160
rect 38204 52096 38220 52160
rect 38284 52156 43740 52160
rect 38284 52100 40165 52156
rect 40221 52100 43055 52156
rect 43111 52100 43740 52156
rect 38284 52096 43740 52100
rect 43804 52096 43820 52160
rect 43884 52096 43900 52160
rect 43964 52096 43980 52160
rect 44044 52096 44060 52160
rect 44124 52096 44140 52160
rect 44204 52096 44220 52160
rect 44284 52156 49740 52160
rect 49804 52156 49820 52160
rect 49884 52156 49900 52160
rect 44284 52100 45945 52156
rect 46001 52100 48892 52156
rect 48948 52100 49740 52156
rect 49810 52100 49820 52156
rect 49890 52100 49900 52156
rect 44284 52096 49740 52100
rect 49804 52096 49820 52100
rect 49884 52096 49900 52100
rect 49964 52096 49980 52160
rect 50044 52096 50060 52160
rect 50124 52096 50140 52160
rect 50204 52096 50220 52160
rect 50284 52156 55740 52160
rect 50284 52100 53048 52156
rect 53104 52100 53206 52156
rect 53262 52100 53562 52156
rect 53618 52100 54880 52156
rect 54936 52100 55473 52156
rect 55529 52100 55740 52156
rect 50284 52096 55740 52100
rect 55804 52096 55820 52160
rect 55884 52096 55900 52160
rect 55964 52096 55980 52160
rect 56044 52096 56060 52160
rect 56124 52096 56140 52160
rect 56204 52096 56220 52160
rect 56284 52156 61740 52160
rect 56284 52100 56619 52156
rect 56675 52100 58055 52156
rect 58111 52100 58135 52156
rect 58191 52100 59298 52156
rect 59354 52100 59456 52156
rect 59512 52100 59764 52156
rect 59820 52100 59910 52156
rect 59966 52100 60046 52156
rect 60102 52100 60126 52156
rect 60182 52100 61740 52156
rect 56284 52096 61740 52100
rect 61804 52096 61820 52160
rect 61884 52096 61900 52160
rect 61964 52096 61980 52160
rect 62044 52096 62060 52160
rect 62124 52096 62140 52160
rect 62204 52096 62220 52160
rect 62284 52156 67740 52160
rect 62284 52100 62418 52156
rect 62474 52100 62498 52156
rect 62554 52100 67740 52156
rect 62284 52096 67740 52100
rect 67804 52096 67820 52160
rect 67884 52096 67900 52160
rect 67964 52096 67980 52160
rect 68044 52096 68060 52160
rect 68124 52096 68140 52160
rect 68204 52096 68220 52160
rect 68284 52156 73740 52160
rect 68284 52100 71864 52156
rect 71920 52100 71944 52156
rect 72000 52100 72024 52156
rect 72080 52100 72104 52156
rect 72160 52100 73740 52156
rect 68284 52096 73740 52100
rect 73804 52096 73820 52160
rect 73884 52096 73900 52160
rect 73964 52096 73980 52160
rect 74044 52096 74060 52160
rect 74124 52096 74140 52160
rect 74204 52096 74220 52160
rect 74284 52096 75028 52160
rect 964 52080 75028 52096
rect 964 52016 1740 52080
rect 1804 52016 1820 52080
rect 1884 52016 1900 52080
rect 1964 52016 1980 52080
rect 2044 52016 2060 52080
rect 2124 52016 2140 52080
rect 2204 52016 2220 52080
rect 2284 52076 7740 52080
rect 2332 52020 2356 52076
rect 2412 52020 5485 52076
rect 5541 52020 7740 52076
rect 2284 52016 7740 52020
rect 7804 52016 7820 52080
rect 7884 52016 7900 52080
rect 7964 52016 7980 52080
rect 8044 52016 8060 52080
rect 8124 52016 8140 52080
rect 8204 52016 8220 52080
rect 8284 52076 13740 52080
rect 8284 52020 8375 52076
rect 8431 52020 11265 52076
rect 11321 52020 13740 52076
rect 8284 52016 13740 52020
rect 13804 52016 13820 52080
rect 13884 52016 13900 52080
rect 13964 52016 13980 52080
rect 14044 52016 14060 52080
rect 14124 52016 14140 52080
rect 14204 52076 14220 52080
rect 14211 52020 14220 52076
rect 14204 52016 14220 52020
rect 14284 52076 19740 52080
rect 14284 52020 17045 52076
rect 17101 52020 19740 52076
rect 14284 52016 19740 52020
rect 19804 52016 19820 52080
rect 19884 52016 19900 52080
rect 19964 52076 19980 52080
rect 19964 52016 19980 52020
rect 20044 52016 20060 52080
rect 20124 52016 20140 52080
rect 20204 52016 20220 52080
rect 20284 52076 25740 52080
rect 20284 52020 22825 52076
rect 22881 52020 25715 52076
rect 20284 52016 25740 52020
rect 25804 52016 25820 52080
rect 25884 52016 25900 52080
rect 25964 52016 25980 52080
rect 26044 52016 26060 52080
rect 26124 52016 26140 52080
rect 26204 52016 26220 52080
rect 26284 52076 31740 52080
rect 26284 52020 28605 52076
rect 28661 52020 31495 52076
rect 31551 52020 31740 52076
rect 26284 52016 31740 52020
rect 31804 52016 31820 52080
rect 31884 52016 31900 52080
rect 31964 52016 31980 52080
rect 32044 52016 32060 52080
rect 32124 52016 32140 52080
rect 32204 52016 32220 52080
rect 32284 52076 37740 52080
rect 32284 52020 34385 52076
rect 34441 52020 37275 52076
rect 37331 52020 37740 52076
rect 32284 52016 37740 52020
rect 37804 52016 37820 52080
rect 37884 52016 37900 52080
rect 37964 52016 37980 52080
rect 38044 52016 38060 52080
rect 38124 52016 38140 52080
rect 38204 52016 38220 52080
rect 38284 52076 43740 52080
rect 38284 52020 40165 52076
rect 40221 52020 43055 52076
rect 43111 52020 43740 52076
rect 38284 52016 43740 52020
rect 43804 52016 43820 52080
rect 43884 52016 43900 52080
rect 43964 52016 43980 52080
rect 44044 52016 44060 52080
rect 44124 52016 44140 52080
rect 44204 52016 44220 52080
rect 44284 52076 49740 52080
rect 49804 52076 49820 52080
rect 49884 52076 49900 52080
rect 44284 52020 45945 52076
rect 46001 52020 48892 52076
rect 48948 52020 49740 52076
rect 49810 52020 49820 52076
rect 49890 52020 49900 52076
rect 44284 52016 49740 52020
rect 49804 52016 49820 52020
rect 49884 52016 49900 52020
rect 49964 52016 49980 52080
rect 50044 52016 50060 52080
rect 50124 52016 50140 52080
rect 50204 52016 50220 52080
rect 50284 52076 55740 52080
rect 50284 52020 53048 52076
rect 53104 52020 53206 52076
rect 53262 52020 53562 52076
rect 53618 52020 54880 52076
rect 54936 52020 55473 52076
rect 55529 52020 55740 52076
rect 50284 52016 55740 52020
rect 55804 52016 55820 52080
rect 55884 52016 55900 52080
rect 55964 52016 55980 52080
rect 56044 52016 56060 52080
rect 56124 52016 56140 52080
rect 56204 52016 56220 52080
rect 56284 52076 61740 52080
rect 56284 52020 56619 52076
rect 56675 52020 58055 52076
rect 58111 52020 58135 52076
rect 58191 52020 59298 52076
rect 59354 52020 59456 52076
rect 59512 52020 59764 52076
rect 59820 52020 59910 52076
rect 59966 52020 60046 52076
rect 60102 52020 60126 52076
rect 60182 52020 61740 52076
rect 56284 52016 61740 52020
rect 61804 52016 61820 52080
rect 61884 52016 61900 52080
rect 61964 52016 61980 52080
rect 62044 52016 62060 52080
rect 62124 52016 62140 52080
rect 62204 52016 62220 52080
rect 62284 52076 67740 52080
rect 62284 52020 62418 52076
rect 62474 52020 62498 52076
rect 62554 52020 67740 52076
rect 62284 52016 67740 52020
rect 67804 52016 67820 52080
rect 67884 52016 67900 52080
rect 67964 52016 67980 52080
rect 68044 52016 68060 52080
rect 68124 52016 68140 52080
rect 68204 52016 68220 52080
rect 68284 52076 73740 52080
rect 68284 52020 71864 52076
rect 71920 52020 71944 52076
rect 72000 52020 72024 52076
rect 72080 52020 72104 52076
rect 72160 52020 73740 52076
rect 68284 52016 73740 52020
rect 73804 52016 73820 52080
rect 73884 52016 73900 52080
rect 73964 52016 73980 52080
rect 74044 52016 74060 52080
rect 74124 52016 74140 52080
rect 74204 52016 74220 52080
rect 74284 52016 75028 52080
rect 964 52000 75028 52016
rect 964 51936 1740 52000
rect 1804 51936 1820 52000
rect 1884 51936 1900 52000
rect 1964 51936 1980 52000
rect 2044 51936 2060 52000
rect 2124 51936 2140 52000
rect 2204 51936 2220 52000
rect 2284 51996 7740 52000
rect 2332 51940 2356 51996
rect 2412 51940 5485 51996
rect 5541 51940 7740 51996
rect 2284 51936 7740 51940
rect 7804 51936 7820 52000
rect 7884 51936 7900 52000
rect 7964 51936 7980 52000
rect 8044 51936 8060 52000
rect 8124 51936 8140 52000
rect 8204 51936 8220 52000
rect 8284 51996 13740 52000
rect 8284 51940 8375 51996
rect 8431 51940 11265 51996
rect 11321 51940 13740 51996
rect 8284 51936 13740 51940
rect 13804 51936 13820 52000
rect 13884 51936 13900 52000
rect 13964 51936 13980 52000
rect 14044 51936 14060 52000
rect 14124 51936 14140 52000
rect 14204 51996 14220 52000
rect 14211 51940 14220 51996
rect 14204 51936 14220 51940
rect 14284 51996 19740 52000
rect 14284 51940 17045 51996
rect 17101 51940 19740 51996
rect 14284 51936 19740 51940
rect 19804 51936 19820 52000
rect 19884 51936 19900 52000
rect 19964 51996 19980 52000
rect 19964 51936 19980 51940
rect 20044 51936 20060 52000
rect 20124 51936 20140 52000
rect 20204 51936 20220 52000
rect 20284 51996 25740 52000
rect 20284 51940 22825 51996
rect 22881 51940 25715 51996
rect 20284 51936 25740 51940
rect 25804 51936 25820 52000
rect 25884 51936 25900 52000
rect 25964 51936 25980 52000
rect 26044 51936 26060 52000
rect 26124 51936 26140 52000
rect 26204 51936 26220 52000
rect 26284 51996 31740 52000
rect 26284 51940 28605 51996
rect 28661 51940 31495 51996
rect 31551 51940 31740 51996
rect 26284 51936 31740 51940
rect 31804 51936 31820 52000
rect 31884 51936 31900 52000
rect 31964 51936 31980 52000
rect 32044 51936 32060 52000
rect 32124 51936 32140 52000
rect 32204 51936 32220 52000
rect 32284 51996 37740 52000
rect 32284 51940 34385 51996
rect 34441 51940 37275 51996
rect 37331 51940 37740 51996
rect 32284 51936 37740 51940
rect 37804 51936 37820 52000
rect 37884 51936 37900 52000
rect 37964 51936 37980 52000
rect 38044 51936 38060 52000
rect 38124 51936 38140 52000
rect 38204 51936 38220 52000
rect 38284 51996 43740 52000
rect 38284 51940 40165 51996
rect 40221 51940 43055 51996
rect 43111 51940 43740 51996
rect 38284 51936 43740 51940
rect 43804 51936 43820 52000
rect 43884 51936 43900 52000
rect 43964 51936 43980 52000
rect 44044 51936 44060 52000
rect 44124 51936 44140 52000
rect 44204 51936 44220 52000
rect 44284 51996 49740 52000
rect 49804 51996 49820 52000
rect 49884 51996 49900 52000
rect 44284 51940 45945 51996
rect 46001 51940 48892 51996
rect 48948 51940 49740 51996
rect 49810 51940 49820 51996
rect 49890 51940 49900 51996
rect 44284 51936 49740 51940
rect 49804 51936 49820 51940
rect 49884 51936 49900 51940
rect 49964 51936 49980 52000
rect 50044 51936 50060 52000
rect 50124 51936 50140 52000
rect 50204 51936 50220 52000
rect 50284 51996 55740 52000
rect 50284 51940 53048 51996
rect 53104 51940 53206 51996
rect 53262 51940 53562 51996
rect 53618 51940 54880 51996
rect 54936 51940 55473 51996
rect 55529 51940 55740 51996
rect 50284 51936 55740 51940
rect 55804 51936 55820 52000
rect 55884 51936 55900 52000
rect 55964 51936 55980 52000
rect 56044 51936 56060 52000
rect 56124 51936 56140 52000
rect 56204 51936 56220 52000
rect 56284 51996 61740 52000
rect 56284 51940 56619 51996
rect 56675 51940 58055 51996
rect 58111 51940 58135 51996
rect 58191 51940 59298 51996
rect 59354 51940 59456 51996
rect 59512 51940 59764 51996
rect 59820 51940 59910 51996
rect 59966 51940 60046 51996
rect 60102 51940 60126 51996
rect 60182 51940 61740 51996
rect 56284 51936 61740 51940
rect 61804 51936 61820 52000
rect 61884 51936 61900 52000
rect 61964 51936 61980 52000
rect 62044 51936 62060 52000
rect 62124 51936 62140 52000
rect 62204 51936 62220 52000
rect 62284 51996 67740 52000
rect 62284 51940 62418 51996
rect 62474 51940 62498 51996
rect 62554 51940 67740 51996
rect 62284 51936 67740 51940
rect 67804 51936 67820 52000
rect 67884 51936 67900 52000
rect 67964 51936 67980 52000
rect 68044 51936 68060 52000
rect 68124 51936 68140 52000
rect 68204 51936 68220 52000
rect 68284 51996 73740 52000
rect 68284 51940 71864 51996
rect 71920 51940 71944 51996
rect 72000 51940 72024 51996
rect 72080 51940 72104 51996
rect 72160 51940 73740 51996
rect 68284 51936 73740 51940
rect 73804 51936 73820 52000
rect 73884 51936 73900 52000
rect 73964 51936 73980 52000
rect 74044 51936 74060 52000
rect 74124 51936 74140 52000
rect 74204 51936 74220 52000
rect 74284 51936 75028 52000
rect 964 51912 75028 51936
rect 65701 47020 65767 47021
rect 65701 47016 65748 47020
rect 65812 47018 65818 47020
rect 65977 47018 66043 47021
rect 66110 47018 66116 47020
rect 65701 46960 65706 47016
rect 65701 46956 65748 46960
rect 65812 46958 65858 47018
rect 65977 47016 66116 47018
rect 65977 46960 65982 47016
rect 66038 46960 66116 47016
rect 65977 46958 66116 46960
rect 65812 46956 65818 46958
rect 65701 46955 65767 46956
rect 65977 46955 66043 46958
rect 66110 46956 66116 46958
rect 66180 46956 66186 47020
rect 964 44592 75028 44616
rect 964 44588 4740 44592
rect 964 44532 2136 44588
rect 2192 44532 4740 44588
rect 964 44528 4740 44532
rect 4804 44528 4820 44592
rect 4884 44528 4900 44592
rect 4964 44528 4980 44592
rect 5044 44528 5060 44592
rect 5124 44528 5140 44592
rect 5204 44528 5220 44592
rect 5284 44588 10740 44592
rect 5284 44532 5632 44588
rect 5688 44532 8522 44588
rect 8578 44532 10740 44588
rect 5284 44528 10740 44532
rect 10804 44528 10820 44592
rect 10884 44528 10900 44592
rect 10964 44528 10980 44592
rect 11044 44528 11060 44592
rect 11124 44528 11140 44592
rect 11204 44528 11220 44592
rect 11284 44588 16740 44592
rect 11284 44532 11412 44588
rect 11468 44532 14302 44588
rect 14358 44532 16740 44588
rect 11284 44528 16740 44532
rect 16804 44528 16820 44592
rect 16884 44528 16900 44592
rect 16964 44528 16980 44592
rect 17044 44528 17060 44592
rect 17124 44528 17140 44592
rect 17204 44588 17220 44592
rect 17284 44588 22740 44592
rect 17284 44532 20082 44588
rect 20138 44532 22740 44588
rect 17204 44528 17220 44532
rect 17284 44528 22740 44532
rect 22804 44528 22820 44592
rect 22884 44528 22900 44592
rect 22964 44588 22980 44592
rect 22964 44532 22972 44588
rect 22964 44528 22980 44532
rect 23044 44528 23060 44592
rect 23124 44528 23140 44592
rect 23204 44528 23220 44592
rect 23284 44588 28740 44592
rect 28804 44588 28820 44592
rect 23284 44532 25862 44588
rect 25918 44532 28740 44588
rect 28808 44532 28820 44588
rect 23284 44528 28740 44532
rect 28804 44528 28820 44532
rect 28884 44528 28900 44592
rect 28964 44528 28980 44592
rect 29044 44528 29060 44592
rect 29124 44528 29140 44592
rect 29204 44528 29220 44592
rect 29284 44588 34740 44592
rect 29284 44532 31642 44588
rect 31698 44532 34532 44588
rect 34588 44532 34740 44588
rect 29284 44528 34740 44532
rect 34804 44528 34820 44592
rect 34884 44528 34900 44592
rect 34964 44528 34980 44592
rect 35044 44528 35060 44592
rect 35124 44528 35140 44592
rect 35204 44528 35220 44592
rect 35284 44588 40740 44592
rect 35284 44532 37422 44588
rect 37478 44532 40312 44588
rect 40368 44532 40740 44588
rect 35284 44528 40740 44532
rect 40804 44528 40820 44592
rect 40884 44528 40900 44592
rect 40964 44528 40980 44592
rect 41044 44528 41060 44592
rect 41124 44528 41140 44592
rect 41204 44528 41220 44592
rect 41284 44588 46740 44592
rect 41284 44532 43202 44588
rect 43258 44532 46092 44588
rect 46148 44532 46740 44588
rect 41284 44528 46740 44532
rect 46804 44528 46820 44592
rect 46884 44528 46900 44592
rect 46964 44528 46980 44592
rect 47044 44528 47060 44592
rect 47124 44528 47140 44592
rect 47204 44528 47220 44592
rect 47284 44588 52740 44592
rect 47284 44532 52329 44588
rect 52385 44532 52740 44588
rect 47284 44528 52740 44532
rect 52804 44528 52820 44592
rect 52884 44528 52900 44592
rect 52964 44528 52980 44592
rect 53044 44528 53060 44592
rect 53124 44528 53140 44592
rect 53204 44528 53220 44592
rect 53284 44588 58740 44592
rect 53284 44532 53730 44588
rect 53786 44532 54642 44588
rect 54698 44532 55032 44588
rect 55088 44532 55748 44588
rect 55804 44532 56326 44588
rect 56382 44532 56771 44588
rect 56827 44532 57075 44588
rect 57131 44532 57917 44588
rect 57973 44532 58441 44588
rect 58497 44532 58740 44588
rect 53284 44528 58740 44532
rect 58804 44528 58820 44592
rect 58884 44528 58900 44592
rect 58964 44528 58980 44592
rect 59044 44528 59060 44592
rect 59124 44528 59140 44592
rect 59204 44528 59220 44592
rect 59284 44588 64740 44592
rect 59284 44532 60418 44588
rect 60474 44532 60576 44588
rect 60632 44532 62620 44588
rect 62676 44532 62700 44588
rect 62756 44532 64740 44588
rect 59284 44528 64740 44532
rect 64804 44528 64820 44592
rect 64884 44528 64900 44592
rect 64964 44528 64980 44592
rect 65044 44528 65060 44592
rect 65124 44528 65140 44592
rect 65204 44528 65220 44592
rect 65284 44528 70740 44592
rect 70804 44528 70820 44592
rect 70884 44528 70900 44592
rect 70964 44528 70980 44592
rect 71044 44528 71060 44592
rect 71124 44528 71140 44592
rect 71204 44528 71220 44592
rect 71284 44588 75028 44592
rect 71284 44532 74216 44588
rect 74272 44532 74296 44588
rect 74352 44532 74376 44588
rect 74432 44532 74456 44588
rect 74512 44532 75028 44588
rect 71284 44528 75028 44532
rect 964 44512 75028 44528
rect 964 44508 4740 44512
rect 964 44452 2136 44508
rect 2192 44452 4740 44508
rect 964 44448 4740 44452
rect 4804 44448 4820 44512
rect 4884 44448 4900 44512
rect 4964 44448 4980 44512
rect 5044 44448 5060 44512
rect 5124 44448 5140 44512
rect 5204 44448 5220 44512
rect 5284 44508 10740 44512
rect 5284 44452 5632 44508
rect 5688 44452 8522 44508
rect 8578 44452 10740 44508
rect 5284 44448 10740 44452
rect 10804 44448 10820 44512
rect 10884 44448 10900 44512
rect 10964 44448 10980 44512
rect 11044 44448 11060 44512
rect 11124 44448 11140 44512
rect 11204 44448 11220 44512
rect 11284 44508 16740 44512
rect 11284 44452 11412 44508
rect 11468 44452 14302 44508
rect 14358 44452 16740 44508
rect 11284 44448 16740 44452
rect 16804 44448 16820 44512
rect 16884 44448 16900 44512
rect 16964 44448 16980 44512
rect 17044 44448 17060 44512
rect 17124 44448 17140 44512
rect 17204 44508 17220 44512
rect 17284 44508 22740 44512
rect 17284 44452 20082 44508
rect 20138 44452 22740 44508
rect 17204 44448 17220 44452
rect 17284 44448 22740 44452
rect 22804 44448 22820 44512
rect 22884 44448 22900 44512
rect 22964 44508 22980 44512
rect 22964 44452 22972 44508
rect 22964 44448 22980 44452
rect 23044 44448 23060 44512
rect 23124 44448 23140 44512
rect 23204 44448 23220 44512
rect 23284 44508 28740 44512
rect 28804 44508 28820 44512
rect 23284 44452 25862 44508
rect 25918 44452 28740 44508
rect 28808 44452 28820 44508
rect 23284 44448 28740 44452
rect 28804 44448 28820 44452
rect 28884 44448 28900 44512
rect 28964 44448 28980 44512
rect 29044 44448 29060 44512
rect 29124 44448 29140 44512
rect 29204 44448 29220 44512
rect 29284 44508 34740 44512
rect 29284 44452 31642 44508
rect 31698 44452 34532 44508
rect 34588 44452 34740 44508
rect 29284 44448 34740 44452
rect 34804 44448 34820 44512
rect 34884 44448 34900 44512
rect 34964 44448 34980 44512
rect 35044 44448 35060 44512
rect 35124 44448 35140 44512
rect 35204 44448 35220 44512
rect 35284 44508 40740 44512
rect 35284 44452 37422 44508
rect 37478 44452 40312 44508
rect 40368 44452 40740 44508
rect 35284 44448 40740 44452
rect 40804 44448 40820 44512
rect 40884 44448 40900 44512
rect 40964 44448 40980 44512
rect 41044 44448 41060 44512
rect 41124 44448 41140 44512
rect 41204 44448 41220 44512
rect 41284 44508 46740 44512
rect 41284 44452 43202 44508
rect 43258 44452 46092 44508
rect 46148 44452 46740 44508
rect 41284 44448 46740 44452
rect 46804 44448 46820 44512
rect 46884 44448 46900 44512
rect 46964 44448 46980 44512
rect 47044 44448 47060 44512
rect 47124 44448 47140 44512
rect 47204 44448 47220 44512
rect 47284 44508 52740 44512
rect 47284 44452 52329 44508
rect 52385 44452 52740 44508
rect 47284 44448 52740 44452
rect 52804 44448 52820 44512
rect 52884 44448 52900 44512
rect 52964 44448 52980 44512
rect 53044 44448 53060 44512
rect 53124 44448 53140 44512
rect 53204 44448 53220 44512
rect 53284 44508 58740 44512
rect 53284 44452 53730 44508
rect 53786 44452 54642 44508
rect 54698 44452 55032 44508
rect 55088 44452 55748 44508
rect 55804 44452 56326 44508
rect 56382 44452 56771 44508
rect 56827 44452 57075 44508
rect 57131 44452 57917 44508
rect 57973 44452 58441 44508
rect 58497 44452 58740 44508
rect 53284 44448 58740 44452
rect 58804 44448 58820 44512
rect 58884 44448 58900 44512
rect 58964 44448 58980 44512
rect 59044 44448 59060 44512
rect 59124 44448 59140 44512
rect 59204 44448 59220 44512
rect 59284 44508 64740 44512
rect 59284 44452 60418 44508
rect 60474 44452 60576 44508
rect 60632 44452 62620 44508
rect 62676 44452 62700 44508
rect 62756 44452 64740 44508
rect 59284 44448 64740 44452
rect 64804 44448 64820 44512
rect 64884 44448 64900 44512
rect 64964 44448 64980 44512
rect 65044 44448 65060 44512
rect 65124 44448 65140 44512
rect 65204 44448 65220 44512
rect 65284 44448 70740 44512
rect 70804 44448 70820 44512
rect 70884 44448 70900 44512
rect 70964 44448 70980 44512
rect 71044 44448 71060 44512
rect 71124 44448 71140 44512
rect 71204 44448 71220 44512
rect 71284 44508 75028 44512
rect 71284 44452 74216 44508
rect 74272 44452 74296 44508
rect 74352 44452 74376 44508
rect 74432 44452 74456 44508
rect 74512 44452 75028 44508
rect 71284 44448 75028 44452
rect 964 44432 75028 44448
rect 964 44428 4740 44432
rect 964 44372 2136 44428
rect 2192 44372 4740 44428
rect 964 44368 4740 44372
rect 4804 44368 4820 44432
rect 4884 44368 4900 44432
rect 4964 44368 4980 44432
rect 5044 44368 5060 44432
rect 5124 44368 5140 44432
rect 5204 44368 5220 44432
rect 5284 44428 10740 44432
rect 5284 44372 5632 44428
rect 5688 44372 8522 44428
rect 8578 44372 10740 44428
rect 5284 44368 10740 44372
rect 10804 44368 10820 44432
rect 10884 44368 10900 44432
rect 10964 44368 10980 44432
rect 11044 44368 11060 44432
rect 11124 44368 11140 44432
rect 11204 44368 11220 44432
rect 11284 44428 16740 44432
rect 11284 44372 11412 44428
rect 11468 44372 14302 44428
rect 14358 44372 16740 44428
rect 11284 44368 16740 44372
rect 16804 44368 16820 44432
rect 16884 44368 16900 44432
rect 16964 44368 16980 44432
rect 17044 44368 17060 44432
rect 17124 44368 17140 44432
rect 17204 44428 17220 44432
rect 17284 44428 22740 44432
rect 17284 44372 20082 44428
rect 20138 44372 22740 44428
rect 17204 44368 17220 44372
rect 17284 44368 22740 44372
rect 22804 44368 22820 44432
rect 22884 44368 22900 44432
rect 22964 44428 22980 44432
rect 22964 44372 22972 44428
rect 22964 44368 22980 44372
rect 23044 44368 23060 44432
rect 23124 44368 23140 44432
rect 23204 44368 23220 44432
rect 23284 44428 28740 44432
rect 28804 44428 28820 44432
rect 23284 44372 25862 44428
rect 25918 44372 28740 44428
rect 28808 44372 28820 44428
rect 23284 44368 28740 44372
rect 28804 44368 28820 44372
rect 28884 44368 28900 44432
rect 28964 44368 28980 44432
rect 29044 44368 29060 44432
rect 29124 44368 29140 44432
rect 29204 44368 29220 44432
rect 29284 44428 34740 44432
rect 29284 44372 31642 44428
rect 31698 44372 34532 44428
rect 34588 44372 34740 44428
rect 29284 44368 34740 44372
rect 34804 44368 34820 44432
rect 34884 44368 34900 44432
rect 34964 44368 34980 44432
rect 35044 44368 35060 44432
rect 35124 44368 35140 44432
rect 35204 44368 35220 44432
rect 35284 44428 40740 44432
rect 35284 44372 37422 44428
rect 37478 44372 40312 44428
rect 40368 44372 40740 44428
rect 35284 44368 40740 44372
rect 40804 44368 40820 44432
rect 40884 44368 40900 44432
rect 40964 44368 40980 44432
rect 41044 44368 41060 44432
rect 41124 44368 41140 44432
rect 41204 44368 41220 44432
rect 41284 44428 46740 44432
rect 41284 44372 43202 44428
rect 43258 44372 46092 44428
rect 46148 44372 46740 44428
rect 41284 44368 46740 44372
rect 46804 44368 46820 44432
rect 46884 44368 46900 44432
rect 46964 44368 46980 44432
rect 47044 44368 47060 44432
rect 47124 44368 47140 44432
rect 47204 44368 47220 44432
rect 47284 44428 52740 44432
rect 47284 44372 52329 44428
rect 52385 44372 52740 44428
rect 47284 44368 52740 44372
rect 52804 44368 52820 44432
rect 52884 44368 52900 44432
rect 52964 44368 52980 44432
rect 53044 44368 53060 44432
rect 53124 44368 53140 44432
rect 53204 44368 53220 44432
rect 53284 44428 58740 44432
rect 53284 44372 53730 44428
rect 53786 44372 54642 44428
rect 54698 44372 55032 44428
rect 55088 44372 55748 44428
rect 55804 44372 56326 44428
rect 56382 44372 56771 44428
rect 56827 44372 57075 44428
rect 57131 44372 57917 44428
rect 57973 44372 58441 44428
rect 58497 44372 58740 44428
rect 53284 44368 58740 44372
rect 58804 44368 58820 44432
rect 58884 44368 58900 44432
rect 58964 44368 58980 44432
rect 59044 44368 59060 44432
rect 59124 44368 59140 44432
rect 59204 44368 59220 44432
rect 59284 44428 64740 44432
rect 59284 44372 60418 44428
rect 60474 44372 60576 44428
rect 60632 44372 62620 44428
rect 62676 44372 62700 44428
rect 62756 44372 64740 44428
rect 59284 44368 64740 44372
rect 64804 44368 64820 44432
rect 64884 44368 64900 44432
rect 64964 44368 64980 44432
rect 65044 44368 65060 44432
rect 65124 44368 65140 44432
rect 65204 44368 65220 44432
rect 65284 44368 70740 44432
rect 70804 44368 70820 44432
rect 70884 44368 70900 44432
rect 70964 44368 70980 44432
rect 71044 44368 71060 44432
rect 71124 44368 71140 44432
rect 71204 44368 71220 44432
rect 71284 44428 75028 44432
rect 71284 44372 74216 44428
rect 74272 44372 74296 44428
rect 74352 44372 74376 44428
rect 74432 44372 74456 44428
rect 74512 44372 75028 44428
rect 71284 44368 75028 44372
rect 964 44352 75028 44368
rect 964 44348 4740 44352
rect 964 44292 2136 44348
rect 2192 44292 4740 44348
rect 964 44288 4740 44292
rect 4804 44288 4820 44352
rect 4884 44288 4900 44352
rect 4964 44288 4980 44352
rect 5044 44288 5060 44352
rect 5124 44288 5140 44352
rect 5204 44288 5220 44352
rect 5284 44348 10740 44352
rect 5284 44292 5632 44348
rect 5688 44292 8522 44348
rect 8578 44292 10740 44348
rect 5284 44288 10740 44292
rect 10804 44288 10820 44352
rect 10884 44288 10900 44352
rect 10964 44288 10980 44352
rect 11044 44288 11060 44352
rect 11124 44288 11140 44352
rect 11204 44288 11220 44352
rect 11284 44348 16740 44352
rect 11284 44292 11412 44348
rect 11468 44292 14302 44348
rect 14358 44292 16740 44348
rect 11284 44288 16740 44292
rect 16804 44288 16820 44352
rect 16884 44288 16900 44352
rect 16964 44288 16980 44352
rect 17044 44288 17060 44352
rect 17124 44288 17140 44352
rect 17204 44348 17220 44352
rect 17284 44348 22740 44352
rect 17284 44292 20082 44348
rect 20138 44292 22740 44348
rect 17204 44288 17220 44292
rect 17284 44288 22740 44292
rect 22804 44288 22820 44352
rect 22884 44288 22900 44352
rect 22964 44348 22980 44352
rect 22964 44292 22972 44348
rect 22964 44288 22980 44292
rect 23044 44288 23060 44352
rect 23124 44288 23140 44352
rect 23204 44288 23220 44352
rect 23284 44348 28740 44352
rect 28804 44348 28820 44352
rect 23284 44292 25862 44348
rect 25918 44292 28740 44348
rect 28808 44292 28820 44348
rect 23284 44288 28740 44292
rect 28804 44288 28820 44292
rect 28884 44288 28900 44352
rect 28964 44288 28980 44352
rect 29044 44288 29060 44352
rect 29124 44288 29140 44352
rect 29204 44288 29220 44352
rect 29284 44348 34740 44352
rect 29284 44292 31642 44348
rect 31698 44292 34532 44348
rect 34588 44292 34740 44348
rect 29284 44288 34740 44292
rect 34804 44288 34820 44352
rect 34884 44288 34900 44352
rect 34964 44288 34980 44352
rect 35044 44288 35060 44352
rect 35124 44288 35140 44352
rect 35204 44288 35220 44352
rect 35284 44348 40740 44352
rect 35284 44292 37422 44348
rect 37478 44292 40312 44348
rect 40368 44292 40740 44348
rect 35284 44288 40740 44292
rect 40804 44288 40820 44352
rect 40884 44288 40900 44352
rect 40964 44288 40980 44352
rect 41044 44288 41060 44352
rect 41124 44288 41140 44352
rect 41204 44288 41220 44352
rect 41284 44348 46740 44352
rect 41284 44292 43202 44348
rect 43258 44292 46092 44348
rect 46148 44292 46740 44348
rect 41284 44288 46740 44292
rect 46804 44288 46820 44352
rect 46884 44288 46900 44352
rect 46964 44288 46980 44352
rect 47044 44288 47060 44352
rect 47124 44288 47140 44352
rect 47204 44288 47220 44352
rect 47284 44348 52740 44352
rect 47284 44292 52329 44348
rect 52385 44292 52740 44348
rect 47284 44288 52740 44292
rect 52804 44288 52820 44352
rect 52884 44288 52900 44352
rect 52964 44288 52980 44352
rect 53044 44288 53060 44352
rect 53124 44288 53140 44352
rect 53204 44288 53220 44352
rect 53284 44348 58740 44352
rect 53284 44292 53730 44348
rect 53786 44292 54642 44348
rect 54698 44292 55032 44348
rect 55088 44292 55748 44348
rect 55804 44292 56326 44348
rect 56382 44292 56771 44348
rect 56827 44292 57075 44348
rect 57131 44292 57917 44348
rect 57973 44292 58441 44348
rect 58497 44292 58740 44348
rect 53284 44288 58740 44292
rect 58804 44288 58820 44352
rect 58884 44288 58900 44352
rect 58964 44288 58980 44352
rect 59044 44288 59060 44352
rect 59124 44288 59140 44352
rect 59204 44288 59220 44352
rect 59284 44348 64740 44352
rect 59284 44292 60418 44348
rect 60474 44292 60576 44348
rect 60632 44292 62620 44348
rect 62676 44292 62700 44348
rect 62756 44292 64740 44348
rect 59284 44288 64740 44292
rect 64804 44288 64820 44352
rect 64884 44288 64900 44352
rect 64964 44288 64980 44352
rect 65044 44288 65060 44352
rect 65124 44288 65140 44352
rect 65204 44288 65220 44352
rect 65284 44288 70740 44352
rect 70804 44288 70820 44352
rect 70884 44288 70900 44352
rect 70964 44288 70980 44352
rect 71044 44288 71060 44352
rect 71124 44288 71140 44352
rect 71204 44288 71220 44352
rect 71284 44348 75028 44352
rect 71284 44292 74216 44348
rect 74272 44292 74296 44348
rect 74352 44292 74376 44348
rect 74432 44292 74456 44348
rect 74512 44292 75028 44348
rect 71284 44288 75028 44292
rect 964 44264 75028 44288
rect 964 42240 75028 42264
rect 964 42176 1740 42240
rect 1804 42176 1820 42240
rect 1884 42176 1900 42240
rect 1964 42176 1980 42240
rect 2044 42176 2060 42240
rect 2124 42176 2140 42240
rect 2204 42176 2220 42240
rect 2284 42236 7740 42240
rect 2332 42180 2356 42236
rect 2412 42180 5485 42236
rect 5541 42180 7740 42236
rect 2284 42176 7740 42180
rect 7804 42176 7820 42240
rect 7884 42176 7900 42240
rect 7964 42176 7980 42240
rect 8044 42176 8060 42240
rect 8124 42176 8140 42240
rect 8204 42176 8220 42240
rect 8284 42236 13740 42240
rect 8284 42180 8375 42236
rect 8431 42180 11265 42236
rect 11321 42180 13740 42236
rect 8284 42176 13740 42180
rect 13804 42176 13820 42240
rect 13884 42176 13900 42240
rect 13964 42176 13980 42240
rect 14044 42176 14060 42240
rect 14124 42176 14140 42240
rect 14204 42236 14220 42240
rect 14211 42180 14220 42236
rect 14204 42176 14220 42180
rect 14284 42236 19740 42240
rect 14284 42180 17045 42236
rect 17101 42180 19740 42236
rect 14284 42176 19740 42180
rect 19804 42176 19820 42240
rect 19884 42176 19900 42240
rect 19964 42236 19980 42240
rect 19964 42176 19980 42180
rect 20044 42176 20060 42240
rect 20124 42176 20140 42240
rect 20204 42176 20220 42240
rect 20284 42236 25740 42240
rect 20284 42180 22825 42236
rect 22881 42180 25715 42236
rect 20284 42176 25740 42180
rect 25804 42176 25820 42240
rect 25884 42176 25900 42240
rect 25964 42176 25980 42240
rect 26044 42176 26060 42240
rect 26124 42176 26140 42240
rect 26204 42176 26220 42240
rect 26284 42236 31740 42240
rect 26284 42180 28605 42236
rect 28661 42180 31495 42236
rect 31551 42180 31740 42236
rect 26284 42176 31740 42180
rect 31804 42176 31820 42240
rect 31884 42176 31900 42240
rect 31964 42176 31980 42240
rect 32044 42176 32060 42240
rect 32124 42176 32140 42240
rect 32204 42176 32220 42240
rect 32284 42236 37740 42240
rect 32284 42180 34385 42236
rect 34441 42180 37275 42236
rect 37331 42180 37740 42236
rect 32284 42176 37740 42180
rect 37804 42176 37820 42240
rect 37884 42176 37900 42240
rect 37964 42176 37980 42240
rect 38044 42176 38060 42240
rect 38124 42176 38140 42240
rect 38204 42176 38220 42240
rect 38284 42236 43740 42240
rect 38284 42180 40165 42236
rect 40221 42180 43055 42236
rect 43111 42180 43740 42236
rect 38284 42176 43740 42180
rect 43804 42176 43820 42240
rect 43884 42176 43900 42240
rect 43964 42176 43980 42240
rect 44044 42176 44060 42240
rect 44124 42176 44140 42240
rect 44204 42176 44220 42240
rect 44284 42236 49740 42240
rect 49804 42236 49820 42240
rect 49884 42236 49900 42240
rect 44284 42180 45945 42236
rect 46001 42180 48892 42236
rect 48948 42180 49740 42236
rect 49810 42180 49820 42236
rect 49890 42180 49900 42236
rect 44284 42176 49740 42180
rect 49804 42176 49820 42180
rect 49884 42176 49900 42180
rect 49964 42176 49980 42240
rect 50044 42176 50060 42240
rect 50124 42176 50140 42240
rect 50204 42176 50220 42240
rect 50284 42236 55740 42240
rect 50284 42180 53048 42236
rect 53104 42180 53206 42236
rect 53262 42180 53562 42236
rect 53618 42180 54880 42236
rect 54936 42180 55473 42236
rect 55529 42180 55740 42236
rect 50284 42176 55740 42180
rect 55804 42176 55820 42240
rect 55884 42176 55900 42240
rect 55964 42176 55980 42240
rect 56044 42176 56060 42240
rect 56124 42176 56140 42240
rect 56204 42176 56220 42240
rect 56284 42236 61740 42240
rect 56284 42180 56619 42236
rect 56675 42180 58055 42236
rect 58111 42180 58135 42236
rect 58191 42180 59298 42236
rect 59354 42180 59456 42236
rect 59512 42180 59764 42236
rect 59820 42180 59910 42236
rect 59966 42180 60046 42236
rect 60102 42180 60126 42236
rect 60182 42180 61740 42236
rect 56284 42176 61740 42180
rect 61804 42176 61820 42240
rect 61884 42176 61900 42240
rect 61964 42176 61980 42240
rect 62044 42176 62060 42240
rect 62124 42176 62140 42240
rect 62204 42176 62220 42240
rect 62284 42236 67740 42240
rect 62284 42180 62418 42236
rect 62474 42180 62498 42236
rect 62554 42180 67740 42236
rect 62284 42176 67740 42180
rect 67804 42176 67820 42240
rect 67884 42176 67900 42240
rect 67964 42176 67980 42240
rect 68044 42176 68060 42240
rect 68124 42176 68140 42240
rect 68204 42176 68220 42240
rect 68284 42236 73740 42240
rect 68284 42180 71864 42236
rect 71920 42180 71944 42236
rect 72000 42180 72024 42236
rect 72080 42180 72104 42236
rect 72160 42180 73740 42236
rect 68284 42176 73740 42180
rect 73804 42176 73820 42240
rect 73884 42176 73900 42240
rect 73964 42176 73980 42240
rect 74044 42176 74060 42240
rect 74124 42176 74140 42240
rect 74204 42176 74220 42240
rect 74284 42176 75028 42240
rect 964 42160 75028 42176
rect 964 42096 1740 42160
rect 1804 42096 1820 42160
rect 1884 42096 1900 42160
rect 1964 42096 1980 42160
rect 2044 42096 2060 42160
rect 2124 42096 2140 42160
rect 2204 42096 2220 42160
rect 2284 42156 7740 42160
rect 2332 42100 2356 42156
rect 2412 42100 5485 42156
rect 5541 42100 7740 42156
rect 2284 42096 7740 42100
rect 7804 42096 7820 42160
rect 7884 42096 7900 42160
rect 7964 42096 7980 42160
rect 8044 42096 8060 42160
rect 8124 42096 8140 42160
rect 8204 42096 8220 42160
rect 8284 42156 13740 42160
rect 8284 42100 8375 42156
rect 8431 42100 11265 42156
rect 11321 42100 13740 42156
rect 8284 42096 13740 42100
rect 13804 42096 13820 42160
rect 13884 42096 13900 42160
rect 13964 42096 13980 42160
rect 14044 42096 14060 42160
rect 14124 42096 14140 42160
rect 14204 42156 14220 42160
rect 14211 42100 14220 42156
rect 14204 42096 14220 42100
rect 14284 42156 19740 42160
rect 14284 42100 17045 42156
rect 17101 42100 19740 42156
rect 14284 42096 19740 42100
rect 19804 42096 19820 42160
rect 19884 42096 19900 42160
rect 19964 42156 19980 42160
rect 19964 42096 19980 42100
rect 20044 42096 20060 42160
rect 20124 42096 20140 42160
rect 20204 42096 20220 42160
rect 20284 42156 25740 42160
rect 20284 42100 22825 42156
rect 22881 42100 25715 42156
rect 20284 42096 25740 42100
rect 25804 42096 25820 42160
rect 25884 42096 25900 42160
rect 25964 42096 25980 42160
rect 26044 42096 26060 42160
rect 26124 42096 26140 42160
rect 26204 42096 26220 42160
rect 26284 42156 31740 42160
rect 26284 42100 28605 42156
rect 28661 42100 31495 42156
rect 31551 42100 31740 42156
rect 26284 42096 31740 42100
rect 31804 42096 31820 42160
rect 31884 42096 31900 42160
rect 31964 42096 31980 42160
rect 32044 42096 32060 42160
rect 32124 42096 32140 42160
rect 32204 42096 32220 42160
rect 32284 42156 37740 42160
rect 32284 42100 34385 42156
rect 34441 42100 37275 42156
rect 37331 42100 37740 42156
rect 32284 42096 37740 42100
rect 37804 42096 37820 42160
rect 37884 42096 37900 42160
rect 37964 42096 37980 42160
rect 38044 42096 38060 42160
rect 38124 42096 38140 42160
rect 38204 42096 38220 42160
rect 38284 42156 43740 42160
rect 38284 42100 40165 42156
rect 40221 42100 43055 42156
rect 43111 42100 43740 42156
rect 38284 42096 43740 42100
rect 43804 42096 43820 42160
rect 43884 42096 43900 42160
rect 43964 42096 43980 42160
rect 44044 42096 44060 42160
rect 44124 42096 44140 42160
rect 44204 42096 44220 42160
rect 44284 42156 49740 42160
rect 49804 42156 49820 42160
rect 49884 42156 49900 42160
rect 44284 42100 45945 42156
rect 46001 42100 48892 42156
rect 48948 42100 49740 42156
rect 49810 42100 49820 42156
rect 49890 42100 49900 42156
rect 44284 42096 49740 42100
rect 49804 42096 49820 42100
rect 49884 42096 49900 42100
rect 49964 42096 49980 42160
rect 50044 42096 50060 42160
rect 50124 42096 50140 42160
rect 50204 42096 50220 42160
rect 50284 42156 55740 42160
rect 50284 42100 53048 42156
rect 53104 42100 53206 42156
rect 53262 42100 53562 42156
rect 53618 42100 54880 42156
rect 54936 42100 55473 42156
rect 55529 42100 55740 42156
rect 50284 42096 55740 42100
rect 55804 42096 55820 42160
rect 55884 42096 55900 42160
rect 55964 42096 55980 42160
rect 56044 42096 56060 42160
rect 56124 42096 56140 42160
rect 56204 42096 56220 42160
rect 56284 42156 61740 42160
rect 56284 42100 56619 42156
rect 56675 42100 58055 42156
rect 58111 42100 58135 42156
rect 58191 42100 59298 42156
rect 59354 42100 59456 42156
rect 59512 42100 59764 42156
rect 59820 42100 59910 42156
rect 59966 42100 60046 42156
rect 60102 42100 60126 42156
rect 60182 42100 61740 42156
rect 56284 42096 61740 42100
rect 61804 42096 61820 42160
rect 61884 42096 61900 42160
rect 61964 42096 61980 42160
rect 62044 42096 62060 42160
rect 62124 42096 62140 42160
rect 62204 42096 62220 42160
rect 62284 42156 67740 42160
rect 62284 42100 62418 42156
rect 62474 42100 62498 42156
rect 62554 42100 67740 42156
rect 62284 42096 67740 42100
rect 67804 42096 67820 42160
rect 67884 42096 67900 42160
rect 67964 42096 67980 42160
rect 68044 42096 68060 42160
rect 68124 42096 68140 42160
rect 68204 42096 68220 42160
rect 68284 42156 73740 42160
rect 68284 42100 71864 42156
rect 71920 42100 71944 42156
rect 72000 42100 72024 42156
rect 72080 42100 72104 42156
rect 72160 42100 73740 42156
rect 68284 42096 73740 42100
rect 73804 42096 73820 42160
rect 73884 42096 73900 42160
rect 73964 42096 73980 42160
rect 74044 42096 74060 42160
rect 74124 42096 74140 42160
rect 74204 42096 74220 42160
rect 74284 42096 75028 42160
rect 964 42080 75028 42096
rect 964 42016 1740 42080
rect 1804 42016 1820 42080
rect 1884 42016 1900 42080
rect 1964 42016 1980 42080
rect 2044 42016 2060 42080
rect 2124 42016 2140 42080
rect 2204 42016 2220 42080
rect 2284 42076 7740 42080
rect 2332 42020 2356 42076
rect 2412 42020 5485 42076
rect 5541 42020 7740 42076
rect 2284 42016 7740 42020
rect 7804 42016 7820 42080
rect 7884 42016 7900 42080
rect 7964 42016 7980 42080
rect 8044 42016 8060 42080
rect 8124 42016 8140 42080
rect 8204 42016 8220 42080
rect 8284 42076 13740 42080
rect 8284 42020 8375 42076
rect 8431 42020 11265 42076
rect 11321 42020 13740 42076
rect 8284 42016 13740 42020
rect 13804 42016 13820 42080
rect 13884 42016 13900 42080
rect 13964 42016 13980 42080
rect 14044 42016 14060 42080
rect 14124 42016 14140 42080
rect 14204 42076 14220 42080
rect 14211 42020 14220 42076
rect 14204 42016 14220 42020
rect 14284 42076 19740 42080
rect 14284 42020 17045 42076
rect 17101 42020 19740 42076
rect 14284 42016 19740 42020
rect 19804 42016 19820 42080
rect 19884 42016 19900 42080
rect 19964 42076 19980 42080
rect 19964 42016 19980 42020
rect 20044 42016 20060 42080
rect 20124 42016 20140 42080
rect 20204 42016 20220 42080
rect 20284 42076 25740 42080
rect 20284 42020 22825 42076
rect 22881 42020 25715 42076
rect 20284 42016 25740 42020
rect 25804 42016 25820 42080
rect 25884 42016 25900 42080
rect 25964 42016 25980 42080
rect 26044 42016 26060 42080
rect 26124 42016 26140 42080
rect 26204 42016 26220 42080
rect 26284 42076 31740 42080
rect 26284 42020 28605 42076
rect 28661 42020 31495 42076
rect 31551 42020 31740 42076
rect 26284 42016 31740 42020
rect 31804 42016 31820 42080
rect 31884 42016 31900 42080
rect 31964 42016 31980 42080
rect 32044 42016 32060 42080
rect 32124 42016 32140 42080
rect 32204 42016 32220 42080
rect 32284 42076 37740 42080
rect 32284 42020 34385 42076
rect 34441 42020 37275 42076
rect 37331 42020 37740 42076
rect 32284 42016 37740 42020
rect 37804 42016 37820 42080
rect 37884 42016 37900 42080
rect 37964 42016 37980 42080
rect 38044 42016 38060 42080
rect 38124 42016 38140 42080
rect 38204 42016 38220 42080
rect 38284 42076 43740 42080
rect 38284 42020 40165 42076
rect 40221 42020 43055 42076
rect 43111 42020 43740 42076
rect 38284 42016 43740 42020
rect 43804 42016 43820 42080
rect 43884 42016 43900 42080
rect 43964 42016 43980 42080
rect 44044 42016 44060 42080
rect 44124 42016 44140 42080
rect 44204 42016 44220 42080
rect 44284 42076 49740 42080
rect 49804 42076 49820 42080
rect 49884 42076 49900 42080
rect 44284 42020 45945 42076
rect 46001 42020 48892 42076
rect 48948 42020 49740 42076
rect 49810 42020 49820 42076
rect 49890 42020 49900 42076
rect 44284 42016 49740 42020
rect 49804 42016 49820 42020
rect 49884 42016 49900 42020
rect 49964 42016 49980 42080
rect 50044 42016 50060 42080
rect 50124 42016 50140 42080
rect 50204 42016 50220 42080
rect 50284 42076 55740 42080
rect 50284 42020 53048 42076
rect 53104 42020 53206 42076
rect 53262 42020 53562 42076
rect 53618 42020 54880 42076
rect 54936 42020 55473 42076
rect 55529 42020 55740 42076
rect 50284 42016 55740 42020
rect 55804 42016 55820 42080
rect 55884 42016 55900 42080
rect 55964 42016 55980 42080
rect 56044 42016 56060 42080
rect 56124 42016 56140 42080
rect 56204 42016 56220 42080
rect 56284 42076 61740 42080
rect 56284 42020 56619 42076
rect 56675 42020 58055 42076
rect 58111 42020 58135 42076
rect 58191 42020 59298 42076
rect 59354 42020 59456 42076
rect 59512 42020 59764 42076
rect 59820 42020 59910 42076
rect 59966 42020 60046 42076
rect 60102 42020 60126 42076
rect 60182 42020 61740 42076
rect 56284 42016 61740 42020
rect 61804 42016 61820 42080
rect 61884 42016 61900 42080
rect 61964 42016 61980 42080
rect 62044 42016 62060 42080
rect 62124 42016 62140 42080
rect 62204 42016 62220 42080
rect 62284 42076 67740 42080
rect 62284 42020 62418 42076
rect 62474 42020 62498 42076
rect 62554 42020 67740 42076
rect 62284 42016 67740 42020
rect 67804 42016 67820 42080
rect 67884 42016 67900 42080
rect 67964 42016 67980 42080
rect 68044 42016 68060 42080
rect 68124 42016 68140 42080
rect 68204 42016 68220 42080
rect 68284 42076 73740 42080
rect 68284 42020 71864 42076
rect 71920 42020 71944 42076
rect 72000 42020 72024 42076
rect 72080 42020 72104 42076
rect 72160 42020 73740 42076
rect 68284 42016 73740 42020
rect 73804 42016 73820 42080
rect 73884 42016 73900 42080
rect 73964 42016 73980 42080
rect 74044 42016 74060 42080
rect 74124 42016 74140 42080
rect 74204 42016 74220 42080
rect 74284 42016 75028 42080
rect 964 42000 75028 42016
rect 964 41936 1740 42000
rect 1804 41936 1820 42000
rect 1884 41936 1900 42000
rect 1964 41936 1980 42000
rect 2044 41936 2060 42000
rect 2124 41936 2140 42000
rect 2204 41936 2220 42000
rect 2284 41996 7740 42000
rect 2332 41940 2356 41996
rect 2412 41940 5485 41996
rect 5541 41940 7740 41996
rect 2284 41936 7740 41940
rect 7804 41936 7820 42000
rect 7884 41936 7900 42000
rect 7964 41936 7980 42000
rect 8044 41936 8060 42000
rect 8124 41936 8140 42000
rect 8204 41936 8220 42000
rect 8284 41996 13740 42000
rect 8284 41940 8375 41996
rect 8431 41940 11265 41996
rect 11321 41940 13740 41996
rect 8284 41936 13740 41940
rect 13804 41936 13820 42000
rect 13884 41936 13900 42000
rect 13964 41936 13980 42000
rect 14044 41936 14060 42000
rect 14124 41936 14140 42000
rect 14204 41996 14220 42000
rect 14211 41940 14220 41996
rect 14204 41936 14220 41940
rect 14284 41996 19740 42000
rect 14284 41940 17045 41996
rect 17101 41940 19740 41996
rect 14284 41936 19740 41940
rect 19804 41936 19820 42000
rect 19884 41936 19900 42000
rect 19964 41996 19980 42000
rect 19964 41936 19980 41940
rect 20044 41936 20060 42000
rect 20124 41936 20140 42000
rect 20204 41936 20220 42000
rect 20284 41996 25740 42000
rect 20284 41940 22825 41996
rect 22881 41940 25715 41996
rect 20284 41936 25740 41940
rect 25804 41936 25820 42000
rect 25884 41936 25900 42000
rect 25964 41936 25980 42000
rect 26044 41936 26060 42000
rect 26124 41936 26140 42000
rect 26204 41936 26220 42000
rect 26284 41996 31740 42000
rect 26284 41940 28605 41996
rect 28661 41940 31495 41996
rect 31551 41940 31740 41996
rect 26284 41936 31740 41940
rect 31804 41936 31820 42000
rect 31884 41936 31900 42000
rect 31964 41936 31980 42000
rect 32044 41936 32060 42000
rect 32124 41936 32140 42000
rect 32204 41936 32220 42000
rect 32284 41996 37740 42000
rect 32284 41940 34385 41996
rect 34441 41940 37275 41996
rect 37331 41940 37740 41996
rect 32284 41936 37740 41940
rect 37804 41936 37820 42000
rect 37884 41936 37900 42000
rect 37964 41936 37980 42000
rect 38044 41936 38060 42000
rect 38124 41936 38140 42000
rect 38204 41936 38220 42000
rect 38284 41996 43740 42000
rect 38284 41940 40165 41996
rect 40221 41940 43055 41996
rect 43111 41940 43740 41996
rect 38284 41936 43740 41940
rect 43804 41936 43820 42000
rect 43884 41936 43900 42000
rect 43964 41936 43980 42000
rect 44044 41936 44060 42000
rect 44124 41936 44140 42000
rect 44204 41936 44220 42000
rect 44284 41996 49740 42000
rect 49804 41996 49820 42000
rect 49884 41996 49900 42000
rect 44284 41940 45945 41996
rect 46001 41940 48892 41996
rect 48948 41940 49740 41996
rect 49810 41940 49820 41996
rect 49890 41940 49900 41996
rect 44284 41936 49740 41940
rect 49804 41936 49820 41940
rect 49884 41936 49900 41940
rect 49964 41936 49980 42000
rect 50044 41936 50060 42000
rect 50124 41936 50140 42000
rect 50204 41936 50220 42000
rect 50284 41996 55740 42000
rect 50284 41940 53048 41996
rect 53104 41940 53206 41996
rect 53262 41940 53562 41996
rect 53618 41940 54880 41996
rect 54936 41940 55473 41996
rect 55529 41940 55740 41996
rect 50284 41936 55740 41940
rect 55804 41936 55820 42000
rect 55884 41936 55900 42000
rect 55964 41936 55980 42000
rect 56044 41936 56060 42000
rect 56124 41936 56140 42000
rect 56204 41936 56220 42000
rect 56284 41996 61740 42000
rect 56284 41940 56619 41996
rect 56675 41940 58055 41996
rect 58111 41940 58135 41996
rect 58191 41940 59298 41996
rect 59354 41940 59456 41996
rect 59512 41940 59764 41996
rect 59820 41940 59910 41996
rect 59966 41940 60046 41996
rect 60102 41940 60126 41996
rect 60182 41940 61740 41996
rect 56284 41936 61740 41940
rect 61804 41936 61820 42000
rect 61884 41936 61900 42000
rect 61964 41936 61980 42000
rect 62044 41936 62060 42000
rect 62124 41936 62140 42000
rect 62204 41936 62220 42000
rect 62284 41996 67740 42000
rect 62284 41940 62418 41996
rect 62474 41940 62498 41996
rect 62554 41940 67740 41996
rect 62284 41936 67740 41940
rect 67804 41936 67820 42000
rect 67884 41936 67900 42000
rect 67964 41936 67980 42000
rect 68044 41936 68060 42000
rect 68124 41936 68140 42000
rect 68204 41936 68220 42000
rect 68284 41996 73740 42000
rect 68284 41940 71864 41996
rect 71920 41940 71944 41996
rect 72000 41940 72024 41996
rect 72080 41940 72104 41996
rect 72160 41940 73740 41996
rect 68284 41936 73740 41940
rect 73804 41936 73820 42000
rect 73884 41936 73900 42000
rect 73964 41936 73980 42000
rect 74044 41936 74060 42000
rect 74124 41936 74140 42000
rect 74204 41936 74220 42000
rect 74284 41936 75028 42000
rect 964 41912 75028 41936
rect 63861 41306 63927 41309
rect 65558 41306 65564 41308
rect 63861 41304 65564 41306
rect 63861 41248 63866 41304
rect 63922 41248 65564 41304
rect 63861 41246 65564 41248
rect 63861 41243 63927 41246
rect 65558 41244 65564 41246
rect 65628 41244 65634 41308
rect 65558 38524 65564 38588
rect 65628 38586 65634 38588
rect 65701 38586 65767 38589
rect 65628 38584 65767 38586
rect 65628 38528 65706 38584
rect 65762 38528 65767 38584
rect 65628 38526 65767 38528
rect 65628 38524 65634 38526
rect 65701 38523 65767 38526
rect 65425 34778 65491 34781
rect 65558 34778 65564 34780
rect 65425 34776 65564 34778
rect 65425 34720 65430 34776
rect 65486 34720 65564 34776
rect 65425 34718 65564 34720
rect 65425 34715 65491 34718
rect 65558 34716 65564 34718
rect 65628 34716 65634 34780
rect 964 34592 75028 34616
rect 964 34588 4740 34592
rect 964 34532 2136 34588
rect 2192 34532 4740 34588
rect 964 34528 4740 34532
rect 4804 34528 4820 34592
rect 4884 34528 4900 34592
rect 4964 34528 4980 34592
rect 5044 34528 5060 34592
rect 5124 34528 5140 34592
rect 5204 34528 5220 34592
rect 5284 34588 10740 34592
rect 5284 34532 5632 34588
rect 5688 34532 8522 34588
rect 8578 34532 10740 34588
rect 5284 34528 10740 34532
rect 10804 34528 10820 34592
rect 10884 34528 10900 34592
rect 10964 34528 10980 34592
rect 11044 34528 11060 34592
rect 11124 34528 11140 34592
rect 11204 34528 11220 34592
rect 11284 34588 16740 34592
rect 11284 34532 11412 34588
rect 11468 34532 14302 34588
rect 14358 34532 16740 34588
rect 11284 34528 16740 34532
rect 16804 34528 16820 34592
rect 16884 34528 16900 34592
rect 16964 34528 16980 34592
rect 17044 34528 17060 34592
rect 17124 34528 17140 34592
rect 17204 34588 17220 34592
rect 17284 34588 22740 34592
rect 17284 34532 20082 34588
rect 20138 34532 22740 34588
rect 17204 34528 17220 34532
rect 17284 34528 22740 34532
rect 22804 34528 22820 34592
rect 22884 34528 22900 34592
rect 22964 34588 22980 34592
rect 22964 34532 22972 34588
rect 22964 34528 22980 34532
rect 23044 34528 23060 34592
rect 23124 34528 23140 34592
rect 23204 34528 23220 34592
rect 23284 34588 28740 34592
rect 28804 34588 28820 34592
rect 23284 34532 25862 34588
rect 25918 34532 28740 34588
rect 28808 34532 28820 34588
rect 23284 34528 28740 34532
rect 28804 34528 28820 34532
rect 28884 34528 28900 34592
rect 28964 34528 28980 34592
rect 29044 34528 29060 34592
rect 29124 34528 29140 34592
rect 29204 34528 29220 34592
rect 29284 34588 34740 34592
rect 29284 34532 31642 34588
rect 31698 34532 34532 34588
rect 34588 34532 34740 34588
rect 29284 34528 34740 34532
rect 34804 34528 34820 34592
rect 34884 34528 34900 34592
rect 34964 34528 34980 34592
rect 35044 34528 35060 34592
rect 35124 34528 35140 34592
rect 35204 34528 35220 34592
rect 35284 34588 40740 34592
rect 35284 34532 37422 34588
rect 37478 34532 40312 34588
rect 40368 34532 40740 34588
rect 35284 34528 40740 34532
rect 40804 34528 40820 34592
rect 40884 34528 40900 34592
rect 40964 34528 40980 34592
rect 41044 34528 41060 34592
rect 41124 34528 41140 34592
rect 41204 34528 41220 34592
rect 41284 34588 46740 34592
rect 41284 34532 43202 34588
rect 43258 34532 46092 34588
rect 46148 34532 46740 34588
rect 41284 34528 46740 34532
rect 46804 34528 46820 34592
rect 46884 34528 46900 34592
rect 46964 34528 46980 34592
rect 47044 34528 47060 34592
rect 47124 34528 47140 34592
rect 47204 34528 47220 34592
rect 47284 34588 52740 34592
rect 47284 34532 49100 34588
rect 49156 34532 52329 34588
rect 52385 34532 52740 34588
rect 47284 34528 52740 34532
rect 52804 34528 52820 34592
rect 52884 34528 52900 34592
rect 52964 34528 52980 34592
rect 53044 34528 53060 34592
rect 53124 34528 53140 34592
rect 53204 34528 53220 34592
rect 53284 34588 58740 34592
rect 53284 34532 53730 34588
rect 53786 34532 53898 34588
rect 53954 34532 54642 34588
rect 54698 34532 55032 34588
rect 55088 34532 55748 34588
rect 55804 34532 56326 34588
rect 56382 34532 56771 34588
rect 56827 34532 57075 34588
rect 57131 34532 57917 34588
rect 57973 34532 58557 34588
rect 58613 34532 58740 34588
rect 53284 34528 58740 34532
rect 58804 34528 58820 34592
rect 58884 34528 58900 34592
rect 58964 34528 58980 34592
rect 59044 34528 59060 34592
rect 59124 34528 59140 34592
rect 59204 34528 59220 34592
rect 59284 34588 64740 34592
rect 59284 34532 60418 34588
rect 60474 34532 60576 34588
rect 60632 34532 62620 34588
rect 62676 34532 62700 34588
rect 62756 34532 64740 34588
rect 59284 34528 64740 34532
rect 64804 34528 64820 34592
rect 64884 34528 64900 34592
rect 64964 34528 64980 34592
rect 65044 34528 65060 34592
rect 65124 34528 65140 34592
rect 65204 34528 65220 34592
rect 65284 34528 70740 34592
rect 70804 34528 70820 34592
rect 70884 34528 70900 34592
rect 70964 34528 70980 34592
rect 71044 34528 71060 34592
rect 71124 34528 71140 34592
rect 71204 34528 71220 34592
rect 71284 34588 75028 34592
rect 71284 34532 74216 34588
rect 74272 34532 74296 34588
rect 74352 34532 74376 34588
rect 74432 34532 74456 34588
rect 74512 34532 75028 34588
rect 71284 34528 75028 34532
rect 964 34512 75028 34528
rect 964 34508 4740 34512
rect 964 34452 2136 34508
rect 2192 34452 4740 34508
rect 964 34448 4740 34452
rect 4804 34448 4820 34512
rect 4884 34448 4900 34512
rect 4964 34448 4980 34512
rect 5044 34448 5060 34512
rect 5124 34448 5140 34512
rect 5204 34448 5220 34512
rect 5284 34508 10740 34512
rect 5284 34452 5632 34508
rect 5688 34452 8522 34508
rect 8578 34452 10740 34508
rect 5284 34448 10740 34452
rect 10804 34448 10820 34512
rect 10884 34448 10900 34512
rect 10964 34448 10980 34512
rect 11044 34448 11060 34512
rect 11124 34448 11140 34512
rect 11204 34448 11220 34512
rect 11284 34508 16740 34512
rect 11284 34452 11412 34508
rect 11468 34452 14302 34508
rect 14358 34452 16740 34508
rect 11284 34448 16740 34452
rect 16804 34448 16820 34512
rect 16884 34448 16900 34512
rect 16964 34448 16980 34512
rect 17044 34448 17060 34512
rect 17124 34448 17140 34512
rect 17204 34508 17220 34512
rect 17284 34508 22740 34512
rect 17284 34452 20082 34508
rect 20138 34452 22740 34508
rect 17204 34448 17220 34452
rect 17284 34448 22740 34452
rect 22804 34448 22820 34512
rect 22884 34448 22900 34512
rect 22964 34508 22980 34512
rect 22964 34452 22972 34508
rect 22964 34448 22980 34452
rect 23044 34448 23060 34512
rect 23124 34448 23140 34512
rect 23204 34448 23220 34512
rect 23284 34508 28740 34512
rect 28804 34508 28820 34512
rect 23284 34452 25862 34508
rect 25918 34452 28740 34508
rect 28808 34452 28820 34508
rect 23284 34448 28740 34452
rect 28804 34448 28820 34452
rect 28884 34448 28900 34512
rect 28964 34448 28980 34512
rect 29044 34448 29060 34512
rect 29124 34448 29140 34512
rect 29204 34448 29220 34512
rect 29284 34508 34740 34512
rect 29284 34452 31642 34508
rect 31698 34452 34532 34508
rect 34588 34452 34740 34508
rect 29284 34448 34740 34452
rect 34804 34448 34820 34512
rect 34884 34448 34900 34512
rect 34964 34448 34980 34512
rect 35044 34448 35060 34512
rect 35124 34448 35140 34512
rect 35204 34448 35220 34512
rect 35284 34508 40740 34512
rect 35284 34452 37422 34508
rect 37478 34452 40312 34508
rect 40368 34452 40740 34508
rect 35284 34448 40740 34452
rect 40804 34448 40820 34512
rect 40884 34448 40900 34512
rect 40964 34448 40980 34512
rect 41044 34448 41060 34512
rect 41124 34448 41140 34512
rect 41204 34448 41220 34512
rect 41284 34508 46740 34512
rect 41284 34452 43202 34508
rect 43258 34452 46092 34508
rect 46148 34452 46740 34508
rect 41284 34448 46740 34452
rect 46804 34448 46820 34512
rect 46884 34448 46900 34512
rect 46964 34448 46980 34512
rect 47044 34448 47060 34512
rect 47124 34448 47140 34512
rect 47204 34448 47220 34512
rect 47284 34508 52740 34512
rect 47284 34452 49100 34508
rect 49156 34452 52329 34508
rect 52385 34452 52740 34508
rect 47284 34448 52740 34452
rect 52804 34448 52820 34512
rect 52884 34448 52900 34512
rect 52964 34448 52980 34512
rect 53044 34448 53060 34512
rect 53124 34448 53140 34512
rect 53204 34448 53220 34512
rect 53284 34508 58740 34512
rect 53284 34452 53730 34508
rect 53786 34452 53898 34508
rect 53954 34452 54642 34508
rect 54698 34452 55032 34508
rect 55088 34452 55748 34508
rect 55804 34452 56326 34508
rect 56382 34452 56771 34508
rect 56827 34452 57075 34508
rect 57131 34452 57917 34508
rect 57973 34452 58557 34508
rect 58613 34452 58740 34508
rect 53284 34448 58740 34452
rect 58804 34448 58820 34512
rect 58884 34448 58900 34512
rect 58964 34448 58980 34512
rect 59044 34448 59060 34512
rect 59124 34448 59140 34512
rect 59204 34448 59220 34512
rect 59284 34508 64740 34512
rect 59284 34452 60418 34508
rect 60474 34452 60576 34508
rect 60632 34452 62620 34508
rect 62676 34452 62700 34508
rect 62756 34452 64740 34508
rect 59284 34448 64740 34452
rect 64804 34448 64820 34512
rect 64884 34448 64900 34512
rect 64964 34448 64980 34512
rect 65044 34448 65060 34512
rect 65124 34448 65140 34512
rect 65204 34448 65220 34512
rect 65284 34448 70740 34512
rect 70804 34448 70820 34512
rect 70884 34448 70900 34512
rect 70964 34448 70980 34512
rect 71044 34448 71060 34512
rect 71124 34448 71140 34512
rect 71204 34448 71220 34512
rect 71284 34508 75028 34512
rect 71284 34452 74216 34508
rect 74272 34452 74296 34508
rect 74352 34452 74376 34508
rect 74432 34452 74456 34508
rect 74512 34452 75028 34508
rect 71284 34448 75028 34452
rect 964 34432 75028 34448
rect 964 34428 4740 34432
rect 964 34372 2136 34428
rect 2192 34372 4740 34428
rect 964 34368 4740 34372
rect 4804 34368 4820 34432
rect 4884 34368 4900 34432
rect 4964 34368 4980 34432
rect 5044 34368 5060 34432
rect 5124 34368 5140 34432
rect 5204 34368 5220 34432
rect 5284 34428 10740 34432
rect 5284 34372 5632 34428
rect 5688 34372 8522 34428
rect 8578 34372 10740 34428
rect 5284 34368 10740 34372
rect 10804 34368 10820 34432
rect 10884 34368 10900 34432
rect 10964 34368 10980 34432
rect 11044 34368 11060 34432
rect 11124 34368 11140 34432
rect 11204 34368 11220 34432
rect 11284 34428 16740 34432
rect 11284 34372 11412 34428
rect 11468 34372 14302 34428
rect 14358 34372 16740 34428
rect 11284 34368 16740 34372
rect 16804 34368 16820 34432
rect 16884 34368 16900 34432
rect 16964 34368 16980 34432
rect 17044 34368 17060 34432
rect 17124 34368 17140 34432
rect 17204 34428 17220 34432
rect 17284 34428 22740 34432
rect 17284 34372 20082 34428
rect 20138 34372 22740 34428
rect 17204 34368 17220 34372
rect 17284 34368 22740 34372
rect 22804 34368 22820 34432
rect 22884 34368 22900 34432
rect 22964 34428 22980 34432
rect 22964 34372 22972 34428
rect 22964 34368 22980 34372
rect 23044 34368 23060 34432
rect 23124 34368 23140 34432
rect 23204 34368 23220 34432
rect 23284 34428 28740 34432
rect 28804 34428 28820 34432
rect 23284 34372 25862 34428
rect 25918 34372 28740 34428
rect 28808 34372 28820 34428
rect 23284 34368 28740 34372
rect 28804 34368 28820 34372
rect 28884 34368 28900 34432
rect 28964 34368 28980 34432
rect 29044 34368 29060 34432
rect 29124 34368 29140 34432
rect 29204 34368 29220 34432
rect 29284 34428 34740 34432
rect 29284 34372 31642 34428
rect 31698 34372 34532 34428
rect 34588 34372 34740 34428
rect 29284 34368 34740 34372
rect 34804 34368 34820 34432
rect 34884 34368 34900 34432
rect 34964 34368 34980 34432
rect 35044 34368 35060 34432
rect 35124 34368 35140 34432
rect 35204 34368 35220 34432
rect 35284 34428 40740 34432
rect 35284 34372 37422 34428
rect 37478 34372 40312 34428
rect 40368 34372 40740 34428
rect 35284 34368 40740 34372
rect 40804 34368 40820 34432
rect 40884 34368 40900 34432
rect 40964 34368 40980 34432
rect 41044 34368 41060 34432
rect 41124 34368 41140 34432
rect 41204 34368 41220 34432
rect 41284 34428 46740 34432
rect 41284 34372 43202 34428
rect 43258 34372 46092 34428
rect 46148 34372 46740 34428
rect 41284 34368 46740 34372
rect 46804 34368 46820 34432
rect 46884 34368 46900 34432
rect 46964 34368 46980 34432
rect 47044 34368 47060 34432
rect 47124 34368 47140 34432
rect 47204 34368 47220 34432
rect 47284 34428 52740 34432
rect 47284 34372 49100 34428
rect 49156 34372 52329 34428
rect 52385 34372 52740 34428
rect 47284 34368 52740 34372
rect 52804 34368 52820 34432
rect 52884 34368 52900 34432
rect 52964 34368 52980 34432
rect 53044 34368 53060 34432
rect 53124 34368 53140 34432
rect 53204 34368 53220 34432
rect 53284 34428 58740 34432
rect 53284 34372 53730 34428
rect 53786 34372 53898 34428
rect 53954 34372 54642 34428
rect 54698 34372 55032 34428
rect 55088 34372 55748 34428
rect 55804 34372 56326 34428
rect 56382 34372 56771 34428
rect 56827 34372 57075 34428
rect 57131 34372 57917 34428
rect 57973 34372 58557 34428
rect 58613 34372 58740 34428
rect 53284 34368 58740 34372
rect 58804 34368 58820 34432
rect 58884 34368 58900 34432
rect 58964 34368 58980 34432
rect 59044 34368 59060 34432
rect 59124 34368 59140 34432
rect 59204 34368 59220 34432
rect 59284 34428 64740 34432
rect 59284 34372 60418 34428
rect 60474 34372 60576 34428
rect 60632 34372 62620 34428
rect 62676 34372 62700 34428
rect 62756 34372 64740 34428
rect 59284 34368 64740 34372
rect 64804 34368 64820 34432
rect 64884 34368 64900 34432
rect 64964 34368 64980 34432
rect 65044 34368 65060 34432
rect 65124 34368 65140 34432
rect 65204 34368 65220 34432
rect 65284 34368 70740 34432
rect 70804 34368 70820 34432
rect 70884 34368 70900 34432
rect 70964 34368 70980 34432
rect 71044 34368 71060 34432
rect 71124 34368 71140 34432
rect 71204 34368 71220 34432
rect 71284 34428 75028 34432
rect 71284 34372 74216 34428
rect 74272 34372 74296 34428
rect 74352 34372 74376 34428
rect 74432 34372 74456 34428
rect 74512 34372 75028 34428
rect 71284 34368 75028 34372
rect 964 34352 75028 34368
rect 964 34348 4740 34352
rect 964 34292 2136 34348
rect 2192 34292 4740 34348
rect 964 34288 4740 34292
rect 4804 34288 4820 34352
rect 4884 34288 4900 34352
rect 4964 34288 4980 34352
rect 5044 34288 5060 34352
rect 5124 34288 5140 34352
rect 5204 34288 5220 34352
rect 5284 34348 10740 34352
rect 5284 34292 5632 34348
rect 5688 34292 8522 34348
rect 8578 34292 10740 34348
rect 5284 34288 10740 34292
rect 10804 34288 10820 34352
rect 10884 34288 10900 34352
rect 10964 34288 10980 34352
rect 11044 34288 11060 34352
rect 11124 34288 11140 34352
rect 11204 34288 11220 34352
rect 11284 34348 16740 34352
rect 11284 34292 11412 34348
rect 11468 34292 14302 34348
rect 14358 34292 16740 34348
rect 11284 34288 16740 34292
rect 16804 34288 16820 34352
rect 16884 34288 16900 34352
rect 16964 34288 16980 34352
rect 17044 34288 17060 34352
rect 17124 34288 17140 34352
rect 17204 34348 17220 34352
rect 17284 34348 22740 34352
rect 17284 34292 20082 34348
rect 20138 34292 22740 34348
rect 17204 34288 17220 34292
rect 17284 34288 22740 34292
rect 22804 34288 22820 34352
rect 22884 34288 22900 34352
rect 22964 34348 22980 34352
rect 22964 34292 22972 34348
rect 22964 34288 22980 34292
rect 23044 34288 23060 34352
rect 23124 34288 23140 34352
rect 23204 34288 23220 34352
rect 23284 34348 28740 34352
rect 28804 34348 28820 34352
rect 23284 34292 25862 34348
rect 25918 34292 28740 34348
rect 28808 34292 28820 34348
rect 23284 34288 28740 34292
rect 28804 34288 28820 34292
rect 28884 34288 28900 34352
rect 28964 34288 28980 34352
rect 29044 34288 29060 34352
rect 29124 34288 29140 34352
rect 29204 34288 29220 34352
rect 29284 34348 34740 34352
rect 29284 34292 31642 34348
rect 31698 34292 34532 34348
rect 34588 34292 34740 34348
rect 29284 34288 34740 34292
rect 34804 34288 34820 34352
rect 34884 34288 34900 34352
rect 34964 34288 34980 34352
rect 35044 34288 35060 34352
rect 35124 34288 35140 34352
rect 35204 34288 35220 34352
rect 35284 34348 40740 34352
rect 35284 34292 37422 34348
rect 37478 34292 40312 34348
rect 40368 34292 40740 34348
rect 35284 34288 40740 34292
rect 40804 34288 40820 34352
rect 40884 34288 40900 34352
rect 40964 34288 40980 34352
rect 41044 34288 41060 34352
rect 41124 34288 41140 34352
rect 41204 34288 41220 34352
rect 41284 34348 46740 34352
rect 41284 34292 43202 34348
rect 43258 34292 46092 34348
rect 46148 34292 46740 34348
rect 41284 34288 46740 34292
rect 46804 34288 46820 34352
rect 46884 34288 46900 34352
rect 46964 34288 46980 34352
rect 47044 34288 47060 34352
rect 47124 34288 47140 34352
rect 47204 34288 47220 34352
rect 47284 34348 52740 34352
rect 47284 34292 49100 34348
rect 49156 34292 52329 34348
rect 52385 34292 52740 34348
rect 47284 34288 52740 34292
rect 52804 34288 52820 34352
rect 52884 34288 52900 34352
rect 52964 34288 52980 34352
rect 53044 34288 53060 34352
rect 53124 34288 53140 34352
rect 53204 34288 53220 34352
rect 53284 34348 58740 34352
rect 53284 34292 53730 34348
rect 53786 34292 53898 34348
rect 53954 34292 54642 34348
rect 54698 34292 55032 34348
rect 55088 34292 55748 34348
rect 55804 34292 56326 34348
rect 56382 34292 56771 34348
rect 56827 34292 57075 34348
rect 57131 34292 57917 34348
rect 57973 34292 58557 34348
rect 58613 34292 58740 34348
rect 53284 34288 58740 34292
rect 58804 34288 58820 34352
rect 58884 34288 58900 34352
rect 58964 34288 58980 34352
rect 59044 34288 59060 34352
rect 59124 34288 59140 34352
rect 59204 34288 59220 34352
rect 59284 34348 64740 34352
rect 59284 34292 60418 34348
rect 60474 34292 60576 34348
rect 60632 34292 62620 34348
rect 62676 34292 62700 34348
rect 62756 34292 64740 34348
rect 59284 34288 64740 34292
rect 64804 34288 64820 34352
rect 64884 34288 64900 34352
rect 64964 34288 64980 34352
rect 65044 34288 65060 34352
rect 65124 34288 65140 34352
rect 65204 34288 65220 34352
rect 65284 34288 70740 34352
rect 70804 34288 70820 34352
rect 70884 34288 70900 34352
rect 70964 34288 70980 34352
rect 71044 34288 71060 34352
rect 71124 34288 71140 34352
rect 71204 34288 71220 34352
rect 71284 34348 75028 34352
rect 71284 34292 74216 34348
rect 74272 34292 74296 34348
rect 74352 34292 74376 34348
rect 74432 34292 74456 34348
rect 74512 34292 75028 34348
rect 71284 34288 75028 34292
rect 964 34264 75028 34288
rect 964 32240 75028 32264
rect 964 32176 1740 32240
rect 1804 32176 1820 32240
rect 1884 32176 1900 32240
rect 1964 32176 1980 32240
rect 2044 32176 2060 32240
rect 2124 32176 2140 32240
rect 2204 32176 2220 32240
rect 2284 32236 7740 32240
rect 2332 32180 2356 32236
rect 2412 32180 5485 32236
rect 5541 32180 7740 32236
rect 2284 32176 7740 32180
rect 7804 32176 7820 32240
rect 7884 32176 7900 32240
rect 7964 32176 7980 32240
rect 8044 32176 8060 32240
rect 8124 32176 8140 32240
rect 8204 32176 8220 32240
rect 8284 32236 13740 32240
rect 8284 32180 8375 32236
rect 8431 32180 11265 32236
rect 11321 32180 13740 32236
rect 8284 32176 13740 32180
rect 13804 32176 13820 32240
rect 13884 32176 13900 32240
rect 13964 32176 13980 32240
rect 14044 32176 14060 32240
rect 14124 32176 14140 32240
rect 14204 32236 14220 32240
rect 14211 32180 14220 32236
rect 14204 32176 14220 32180
rect 14284 32236 19740 32240
rect 14284 32180 17045 32236
rect 17101 32180 19740 32236
rect 14284 32176 19740 32180
rect 19804 32176 19820 32240
rect 19884 32176 19900 32240
rect 19964 32236 19980 32240
rect 19964 32176 19980 32180
rect 20044 32176 20060 32240
rect 20124 32176 20140 32240
rect 20204 32176 20220 32240
rect 20284 32236 25740 32240
rect 20284 32180 22825 32236
rect 22881 32180 25715 32236
rect 20284 32176 25740 32180
rect 25804 32176 25820 32240
rect 25884 32176 25900 32240
rect 25964 32176 25980 32240
rect 26044 32176 26060 32240
rect 26124 32176 26140 32240
rect 26204 32176 26220 32240
rect 26284 32236 31740 32240
rect 26284 32180 28605 32236
rect 28661 32180 31495 32236
rect 31551 32180 31740 32236
rect 26284 32176 31740 32180
rect 31804 32176 31820 32240
rect 31884 32176 31900 32240
rect 31964 32176 31980 32240
rect 32044 32176 32060 32240
rect 32124 32176 32140 32240
rect 32204 32176 32220 32240
rect 32284 32236 37740 32240
rect 32284 32180 34385 32236
rect 34441 32180 37275 32236
rect 37331 32180 37740 32236
rect 32284 32176 37740 32180
rect 37804 32176 37820 32240
rect 37884 32176 37900 32240
rect 37964 32176 37980 32240
rect 38044 32176 38060 32240
rect 38124 32176 38140 32240
rect 38204 32176 38220 32240
rect 38284 32236 43740 32240
rect 38284 32180 40165 32236
rect 40221 32180 43055 32236
rect 43111 32180 43740 32236
rect 38284 32176 43740 32180
rect 43804 32176 43820 32240
rect 43884 32176 43900 32240
rect 43964 32176 43980 32240
rect 44044 32176 44060 32240
rect 44124 32176 44140 32240
rect 44204 32176 44220 32240
rect 44284 32236 49740 32240
rect 49804 32236 49820 32240
rect 49884 32236 49900 32240
rect 44284 32180 45945 32236
rect 46001 32180 48892 32236
rect 48948 32180 49740 32236
rect 49810 32180 49820 32236
rect 49890 32180 49900 32236
rect 44284 32176 49740 32180
rect 49804 32176 49820 32180
rect 49884 32176 49900 32180
rect 49964 32176 49980 32240
rect 50044 32176 50060 32240
rect 50124 32176 50140 32240
rect 50204 32176 50220 32240
rect 50284 32236 55740 32240
rect 50284 32180 53048 32236
rect 53104 32180 53206 32236
rect 53262 32180 53562 32236
rect 53618 32180 54880 32236
rect 54936 32180 55473 32236
rect 55529 32180 55740 32236
rect 50284 32176 55740 32180
rect 55804 32176 55820 32240
rect 55884 32176 55900 32240
rect 55964 32176 55980 32240
rect 56044 32176 56060 32240
rect 56124 32176 56140 32240
rect 56204 32176 56220 32240
rect 56284 32236 61740 32240
rect 56284 32180 56619 32236
rect 56675 32180 58055 32236
rect 58111 32180 58135 32236
rect 58191 32180 59298 32236
rect 59354 32180 59456 32236
rect 59512 32180 59764 32236
rect 59820 32180 59910 32236
rect 59966 32180 60046 32236
rect 60102 32180 60126 32236
rect 60182 32180 61740 32236
rect 56284 32176 61740 32180
rect 61804 32176 61820 32240
rect 61884 32176 61900 32240
rect 61964 32176 61980 32240
rect 62044 32176 62060 32240
rect 62124 32176 62140 32240
rect 62204 32176 62220 32240
rect 62284 32236 67740 32240
rect 62284 32180 62418 32236
rect 62474 32180 62498 32236
rect 62554 32180 67740 32236
rect 62284 32176 67740 32180
rect 67804 32176 67820 32240
rect 67884 32176 67900 32240
rect 67964 32176 67980 32240
rect 68044 32176 68060 32240
rect 68124 32176 68140 32240
rect 68204 32176 68220 32240
rect 68284 32236 73740 32240
rect 68284 32180 71864 32236
rect 71920 32180 71944 32236
rect 72000 32180 72024 32236
rect 72080 32180 72104 32236
rect 72160 32180 73740 32236
rect 68284 32176 73740 32180
rect 73804 32176 73820 32240
rect 73884 32176 73900 32240
rect 73964 32176 73980 32240
rect 74044 32176 74060 32240
rect 74124 32176 74140 32240
rect 74204 32176 74220 32240
rect 74284 32176 75028 32240
rect 964 32160 75028 32176
rect 964 32096 1740 32160
rect 1804 32096 1820 32160
rect 1884 32096 1900 32160
rect 1964 32096 1980 32160
rect 2044 32096 2060 32160
rect 2124 32096 2140 32160
rect 2204 32096 2220 32160
rect 2284 32156 7740 32160
rect 2332 32100 2356 32156
rect 2412 32100 5485 32156
rect 5541 32100 7740 32156
rect 2284 32096 7740 32100
rect 7804 32096 7820 32160
rect 7884 32096 7900 32160
rect 7964 32096 7980 32160
rect 8044 32096 8060 32160
rect 8124 32096 8140 32160
rect 8204 32096 8220 32160
rect 8284 32156 13740 32160
rect 8284 32100 8375 32156
rect 8431 32100 11265 32156
rect 11321 32100 13740 32156
rect 8284 32096 13740 32100
rect 13804 32096 13820 32160
rect 13884 32096 13900 32160
rect 13964 32096 13980 32160
rect 14044 32096 14060 32160
rect 14124 32096 14140 32160
rect 14204 32156 14220 32160
rect 14211 32100 14220 32156
rect 14204 32096 14220 32100
rect 14284 32156 19740 32160
rect 14284 32100 17045 32156
rect 17101 32100 19740 32156
rect 14284 32096 19740 32100
rect 19804 32096 19820 32160
rect 19884 32096 19900 32160
rect 19964 32156 19980 32160
rect 19964 32096 19980 32100
rect 20044 32096 20060 32160
rect 20124 32096 20140 32160
rect 20204 32096 20220 32160
rect 20284 32156 25740 32160
rect 20284 32100 22825 32156
rect 22881 32100 25715 32156
rect 20284 32096 25740 32100
rect 25804 32096 25820 32160
rect 25884 32096 25900 32160
rect 25964 32096 25980 32160
rect 26044 32096 26060 32160
rect 26124 32096 26140 32160
rect 26204 32096 26220 32160
rect 26284 32156 31740 32160
rect 26284 32100 28605 32156
rect 28661 32100 31495 32156
rect 31551 32100 31740 32156
rect 26284 32096 31740 32100
rect 31804 32096 31820 32160
rect 31884 32096 31900 32160
rect 31964 32096 31980 32160
rect 32044 32096 32060 32160
rect 32124 32096 32140 32160
rect 32204 32096 32220 32160
rect 32284 32156 37740 32160
rect 32284 32100 34385 32156
rect 34441 32100 37275 32156
rect 37331 32100 37740 32156
rect 32284 32096 37740 32100
rect 37804 32096 37820 32160
rect 37884 32096 37900 32160
rect 37964 32096 37980 32160
rect 38044 32096 38060 32160
rect 38124 32096 38140 32160
rect 38204 32096 38220 32160
rect 38284 32156 43740 32160
rect 38284 32100 40165 32156
rect 40221 32100 43055 32156
rect 43111 32100 43740 32156
rect 38284 32096 43740 32100
rect 43804 32096 43820 32160
rect 43884 32096 43900 32160
rect 43964 32096 43980 32160
rect 44044 32096 44060 32160
rect 44124 32096 44140 32160
rect 44204 32096 44220 32160
rect 44284 32156 49740 32160
rect 49804 32156 49820 32160
rect 49884 32156 49900 32160
rect 44284 32100 45945 32156
rect 46001 32100 48892 32156
rect 48948 32100 49740 32156
rect 49810 32100 49820 32156
rect 49890 32100 49900 32156
rect 44284 32096 49740 32100
rect 49804 32096 49820 32100
rect 49884 32096 49900 32100
rect 49964 32096 49980 32160
rect 50044 32096 50060 32160
rect 50124 32096 50140 32160
rect 50204 32096 50220 32160
rect 50284 32156 55740 32160
rect 50284 32100 53048 32156
rect 53104 32100 53206 32156
rect 53262 32100 53562 32156
rect 53618 32100 54880 32156
rect 54936 32100 55473 32156
rect 55529 32100 55740 32156
rect 50284 32096 55740 32100
rect 55804 32096 55820 32160
rect 55884 32096 55900 32160
rect 55964 32096 55980 32160
rect 56044 32096 56060 32160
rect 56124 32096 56140 32160
rect 56204 32096 56220 32160
rect 56284 32156 61740 32160
rect 56284 32100 56619 32156
rect 56675 32100 58055 32156
rect 58111 32100 58135 32156
rect 58191 32100 59298 32156
rect 59354 32100 59456 32156
rect 59512 32100 59764 32156
rect 59820 32100 59910 32156
rect 59966 32100 60046 32156
rect 60102 32100 60126 32156
rect 60182 32100 61740 32156
rect 56284 32096 61740 32100
rect 61804 32096 61820 32160
rect 61884 32096 61900 32160
rect 61964 32096 61980 32160
rect 62044 32096 62060 32160
rect 62124 32096 62140 32160
rect 62204 32096 62220 32160
rect 62284 32156 67740 32160
rect 62284 32100 62418 32156
rect 62474 32100 62498 32156
rect 62554 32100 67740 32156
rect 62284 32096 67740 32100
rect 67804 32096 67820 32160
rect 67884 32096 67900 32160
rect 67964 32096 67980 32160
rect 68044 32096 68060 32160
rect 68124 32096 68140 32160
rect 68204 32096 68220 32160
rect 68284 32156 73740 32160
rect 68284 32100 71864 32156
rect 71920 32100 71944 32156
rect 72000 32100 72024 32156
rect 72080 32100 72104 32156
rect 72160 32100 73740 32156
rect 68284 32096 73740 32100
rect 73804 32096 73820 32160
rect 73884 32096 73900 32160
rect 73964 32096 73980 32160
rect 74044 32096 74060 32160
rect 74124 32096 74140 32160
rect 74204 32096 74220 32160
rect 74284 32096 75028 32160
rect 964 32080 75028 32096
rect 964 32016 1740 32080
rect 1804 32016 1820 32080
rect 1884 32016 1900 32080
rect 1964 32016 1980 32080
rect 2044 32016 2060 32080
rect 2124 32016 2140 32080
rect 2204 32016 2220 32080
rect 2284 32076 7740 32080
rect 2332 32020 2356 32076
rect 2412 32020 5485 32076
rect 5541 32020 7740 32076
rect 2284 32016 7740 32020
rect 7804 32016 7820 32080
rect 7884 32016 7900 32080
rect 7964 32016 7980 32080
rect 8044 32016 8060 32080
rect 8124 32016 8140 32080
rect 8204 32016 8220 32080
rect 8284 32076 13740 32080
rect 8284 32020 8375 32076
rect 8431 32020 11265 32076
rect 11321 32020 13740 32076
rect 8284 32016 13740 32020
rect 13804 32016 13820 32080
rect 13884 32016 13900 32080
rect 13964 32016 13980 32080
rect 14044 32016 14060 32080
rect 14124 32016 14140 32080
rect 14204 32076 14220 32080
rect 14211 32020 14220 32076
rect 14204 32016 14220 32020
rect 14284 32076 19740 32080
rect 14284 32020 17045 32076
rect 17101 32020 19740 32076
rect 14284 32016 19740 32020
rect 19804 32016 19820 32080
rect 19884 32016 19900 32080
rect 19964 32076 19980 32080
rect 19964 32016 19980 32020
rect 20044 32016 20060 32080
rect 20124 32016 20140 32080
rect 20204 32016 20220 32080
rect 20284 32076 25740 32080
rect 20284 32020 22825 32076
rect 22881 32020 25715 32076
rect 20284 32016 25740 32020
rect 25804 32016 25820 32080
rect 25884 32016 25900 32080
rect 25964 32016 25980 32080
rect 26044 32016 26060 32080
rect 26124 32016 26140 32080
rect 26204 32016 26220 32080
rect 26284 32076 31740 32080
rect 26284 32020 28605 32076
rect 28661 32020 31495 32076
rect 31551 32020 31740 32076
rect 26284 32016 31740 32020
rect 31804 32016 31820 32080
rect 31884 32016 31900 32080
rect 31964 32016 31980 32080
rect 32044 32016 32060 32080
rect 32124 32016 32140 32080
rect 32204 32016 32220 32080
rect 32284 32076 37740 32080
rect 32284 32020 34385 32076
rect 34441 32020 37275 32076
rect 37331 32020 37740 32076
rect 32284 32016 37740 32020
rect 37804 32016 37820 32080
rect 37884 32016 37900 32080
rect 37964 32016 37980 32080
rect 38044 32016 38060 32080
rect 38124 32016 38140 32080
rect 38204 32016 38220 32080
rect 38284 32076 43740 32080
rect 38284 32020 40165 32076
rect 40221 32020 43055 32076
rect 43111 32020 43740 32076
rect 38284 32016 43740 32020
rect 43804 32016 43820 32080
rect 43884 32016 43900 32080
rect 43964 32016 43980 32080
rect 44044 32016 44060 32080
rect 44124 32016 44140 32080
rect 44204 32016 44220 32080
rect 44284 32076 49740 32080
rect 49804 32076 49820 32080
rect 49884 32076 49900 32080
rect 44284 32020 45945 32076
rect 46001 32020 48892 32076
rect 48948 32020 49740 32076
rect 49810 32020 49820 32076
rect 49890 32020 49900 32076
rect 44284 32016 49740 32020
rect 49804 32016 49820 32020
rect 49884 32016 49900 32020
rect 49964 32016 49980 32080
rect 50044 32016 50060 32080
rect 50124 32016 50140 32080
rect 50204 32016 50220 32080
rect 50284 32076 55740 32080
rect 50284 32020 53048 32076
rect 53104 32020 53206 32076
rect 53262 32020 53562 32076
rect 53618 32020 54880 32076
rect 54936 32020 55473 32076
rect 55529 32020 55740 32076
rect 50284 32016 55740 32020
rect 55804 32016 55820 32080
rect 55884 32016 55900 32080
rect 55964 32016 55980 32080
rect 56044 32016 56060 32080
rect 56124 32016 56140 32080
rect 56204 32016 56220 32080
rect 56284 32076 61740 32080
rect 56284 32020 56619 32076
rect 56675 32020 58055 32076
rect 58111 32020 58135 32076
rect 58191 32020 59298 32076
rect 59354 32020 59456 32076
rect 59512 32020 59764 32076
rect 59820 32020 59910 32076
rect 59966 32020 60046 32076
rect 60102 32020 60126 32076
rect 60182 32020 61740 32076
rect 56284 32016 61740 32020
rect 61804 32016 61820 32080
rect 61884 32016 61900 32080
rect 61964 32016 61980 32080
rect 62044 32016 62060 32080
rect 62124 32016 62140 32080
rect 62204 32016 62220 32080
rect 62284 32076 67740 32080
rect 62284 32020 62418 32076
rect 62474 32020 62498 32076
rect 62554 32020 67740 32076
rect 62284 32016 67740 32020
rect 67804 32016 67820 32080
rect 67884 32016 67900 32080
rect 67964 32016 67980 32080
rect 68044 32016 68060 32080
rect 68124 32016 68140 32080
rect 68204 32016 68220 32080
rect 68284 32076 73740 32080
rect 68284 32020 71864 32076
rect 71920 32020 71944 32076
rect 72000 32020 72024 32076
rect 72080 32020 72104 32076
rect 72160 32020 73740 32076
rect 68284 32016 73740 32020
rect 73804 32016 73820 32080
rect 73884 32016 73900 32080
rect 73964 32016 73980 32080
rect 74044 32016 74060 32080
rect 74124 32016 74140 32080
rect 74204 32016 74220 32080
rect 74284 32016 75028 32080
rect 964 32000 75028 32016
rect 964 31936 1740 32000
rect 1804 31936 1820 32000
rect 1884 31936 1900 32000
rect 1964 31936 1980 32000
rect 2044 31936 2060 32000
rect 2124 31936 2140 32000
rect 2204 31936 2220 32000
rect 2284 31996 7740 32000
rect 2332 31940 2356 31996
rect 2412 31940 5485 31996
rect 5541 31940 7740 31996
rect 2284 31936 7740 31940
rect 7804 31936 7820 32000
rect 7884 31936 7900 32000
rect 7964 31936 7980 32000
rect 8044 31936 8060 32000
rect 8124 31936 8140 32000
rect 8204 31936 8220 32000
rect 8284 31996 13740 32000
rect 8284 31940 8375 31996
rect 8431 31940 11265 31996
rect 11321 31940 13740 31996
rect 8284 31936 13740 31940
rect 13804 31936 13820 32000
rect 13884 31936 13900 32000
rect 13964 31936 13980 32000
rect 14044 31936 14060 32000
rect 14124 31936 14140 32000
rect 14204 31996 14220 32000
rect 14211 31940 14220 31996
rect 14204 31936 14220 31940
rect 14284 31996 19740 32000
rect 14284 31940 17045 31996
rect 17101 31940 19740 31996
rect 14284 31936 19740 31940
rect 19804 31936 19820 32000
rect 19884 31936 19900 32000
rect 19964 31996 19980 32000
rect 19964 31936 19980 31940
rect 20044 31936 20060 32000
rect 20124 31936 20140 32000
rect 20204 31936 20220 32000
rect 20284 31996 25740 32000
rect 20284 31940 22825 31996
rect 22881 31940 25715 31996
rect 20284 31936 25740 31940
rect 25804 31936 25820 32000
rect 25884 31936 25900 32000
rect 25964 31936 25980 32000
rect 26044 31936 26060 32000
rect 26124 31936 26140 32000
rect 26204 31936 26220 32000
rect 26284 31996 31740 32000
rect 26284 31940 28605 31996
rect 28661 31940 31495 31996
rect 31551 31940 31740 31996
rect 26284 31936 31740 31940
rect 31804 31936 31820 32000
rect 31884 31936 31900 32000
rect 31964 31936 31980 32000
rect 32044 31936 32060 32000
rect 32124 31936 32140 32000
rect 32204 31936 32220 32000
rect 32284 31996 37740 32000
rect 32284 31940 34385 31996
rect 34441 31940 37275 31996
rect 37331 31940 37740 31996
rect 32284 31936 37740 31940
rect 37804 31936 37820 32000
rect 37884 31936 37900 32000
rect 37964 31936 37980 32000
rect 38044 31936 38060 32000
rect 38124 31936 38140 32000
rect 38204 31936 38220 32000
rect 38284 31996 43740 32000
rect 38284 31940 40165 31996
rect 40221 31940 43055 31996
rect 43111 31940 43740 31996
rect 38284 31936 43740 31940
rect 43804 31936 43820 32000
rect 43884 31936 43900 32000
rect 43964 31936 43980 32000
rect 44044 31936 44060 32000
rect 44124 31936 44140 32000
rect 44204 31936 44220 32000
rect 44284 31996 49740 32000
rect 49804 31996 49820 32000
rect 49884 31996 49900 32000
rect 44284 31940 45945 31996
rect 46001 31940 48892 31996
rect 48948 31940 49740 31996
rect 49810 31940 49820 31996
rect 49890 31940 49900 31996
rect 44284 31936 49740 31940
rect 49804 31936 49820 31940
rect 49884 31936 49900 31940
rect 49964 31936 49980 32000
rect 50044 31936 50060 32000
rect 50124 31936 50140 32000
rect 50204 31936 50220 32000
rect 50284 31996 55740 32000
rect 50284 31940 53048 31996
rect 53104 31940 53206 31996
rect 53262 31940 53562 31996
rect 53618 31940 54880 31996
rect 54936 31940 55473 31996
rect 55529 31940 55740 31996
rect 50284 31936 55740 31940
rect 55804 31936 55820 32000
rect 55884 31936 55900 32000
rect 55964 31936 55980 32000
rect 56044 31936 56060 32000
rect 56124 31936 56140 32000
rect 56204 31936 56220 32000
rect 56284 31996 61740 32000
rect 56284 31940 56619 31996
rect 56675 31940 58055 31996
rect 58111 31940 58135 31996
rect 58191 31940 59298 31996
rect 59354 31940 59456 31996
rect 59512 31940 59764 31996
rect 59820 31940 59910 31996
rect 59966 31940 60046 31996
rect 60102 31940 60126 31996
rect 60182 31940 61740 31996
rect 56284 31936 61740 31940
rect 61804 31936 61820 32000
rect 61884 31936 61900 32000
rect 61964 31936 61980 32000
rect 62044 31936 62060 32000
rect 62124 31936 62140 32000
rect 62204 31936 62220 32000
rect 62284 31996 67740 32000
rect 62284 31940 62418 31996
rect 62474 31940 62498 31996
rect 62554 31940 67740 31996
rect 62284 31936 67740 31940
rect 67804 31936 67820 32000
rect 67884 31936 67900 32000
rect 67964 31936 67980 32000
rect 68044 31936 68060 32000
rect 68124 31936 68140 32000
rect 68204 31936 68220 32000
rect 68284 31996 73740 32000
rect 68284 31940 71864 31996
rect 71920 31940 71944 31996
rect 72000 31940 72024 31996
rect 72080 31940 72104 31996
rect 72160 31940 73740 31996
rect 68284 31936 73740 31940
rect 73804 31936 73820 32000
rect 73884 31936 73900 32000
rect 73964 31936 73980 32000
rect 74044 31936 74060 32000
rect 74124 31936 74140 32000
rect 74204 31936 74220 32000
rect 74284 31936 75028 32000
rect 964 31912 75028 31936
rect 964 24592 75028 24616
rect 964 24588 4740 24592
rect 964 24532 2136 24588
rect 2192 24532 4740 24588
rect 964 24528 4740 24532
rect 4804 24528 4820 24592
rect 4884 24528 4900 24592
rect 4964 24528 4980 24592
rect 5044 24528 5060 24592
rect 5124 24528 5140 24592
rect 5204 24528 5220 24592
rect 5284 24588 10740 24592
rect 5284 24532 5632 24588
rect 5688 24532 8522 24588
rect 8578 24532 10740 24588
rect 5284 24528 10740 24532
rect 10804 24528 10820 24592
rect 10884 24528 10900 24592
rect 10964 24528 10980 24592
rect 11044 24528 11060 24592
rect 11124 24528 11140 24592
rect 11204 24528 11220 24592
rect 11284 24588 16740 24592
rect 11284 24532 11412 24588
rect 11468 24532 14302 24588
rect 14358 24532 16740 24588
rect 11284 24528 16740 24532
rect 16804 24528 16820 24592
rect 16884 24528 16900 24592
rect 16964 24528 16980 24592
rect 17044 24528 17060 24592
rect 17124 24528 17140 24592
rect 17204 24588 17220 24592
rect 17284 24588 22740 24592
rect 17284 24532 20082 24588
rect 20138 24532 22740 24588
rect 17204 24528 17220 24532
rect 17284 24528 22740 24532
rect 22804 24528 22820 24592
rect 22884 24528 22900 24592
rect 22964 24588 22980 24592
rect 22964 24532 22972 24588
rect 22964 24528 22980 24532
rect 23044 24528 23060 24592
rect 23124 24528 23140 24592
rect 23204 24528 23220 24592
rect 23284 24588 28740 24592
rect 28804 24588 28820 24592
rect 23284 24532 25862 24588
rect 25918 24532 28740 24588
rect 28808 24532 28820 24588
rect 23284 24528 28740 24532
rect 28804 24528 28820 24532
rect 28884 24528 28900 24592
rect 28964 24528 28980 24592
rect 29044 24528 29060 24592
rect 29124 24528 29140 24592
rect 29204 24528 29220 24592
rect 29284 24588 34740 24592
rect 29284 24532 31642 24588
rect 31698 24532 34532 24588
rect 34588 24532 34740 24588
rect 29284 24528 34740 24532
rect 34804 24528 34820 24592
rect 34884 24528 34900 24592
rect 34964 24528 34980 24592
rect 35044 24528 35060 24592
rect 35124 24528 35140 24592
rect 35204 24528 35220 24592
rect 35284 24588 40740 24592
rect 35284 24532 37422 24588
rect 37478 24532 40312 24588
rect 40368 24532 40740 24588
rect 35284 24528 40740 24532
rect 40804 24528 40820 24592
rect 40884 24528 40900 24592
rect 40964 24528 40980 24592
rect 41044 24528 41060 24592
rect 41124 24528 41140 24592
rect 41204 24528 41220 24592
rect 41284 24588 46740 24592
rect 41284 24532 43202 24588
rect 43258 24532 46092 24588
rect 46148 24532 46740 24588
rect 41284 24528 46740 24532
rect 46804 24528 46820 24592
rect 46884 24528 46900 24592
rect 46964 24528 46980 24592
rect 47044 24528 47060 24592
rect 47124 24528 47140 24592
rect 47204 24528 47220 24592
rect 47284 24588 52740 24592
rect 47284 24532 49100 24588
rect 49156 24532 52329 24588
rect 52385 24532 52740 24588
rect 47284 24528 52740 24532
rect 52804 24528 52820 24592
rect 52884 24528 52900 24592
rect 52964 24528 52980 24592
rect 53044 24528 53060 24592
rect 53124 24528 53140 24592
rect 53204 24528 53220 24592
rect 53284 24588 58740 24592
rect 53284 24532 53730 24588
rect 53786 24532 53898 24588
rect 53954 24532 54642 24588
rect 54698 24532 55032 24588
rect 55088 24532 55748 24588
rect 55804 24532 56326 24588
rect 56382 24532 56771 24588
rect 56827 24532 57075 24588
rect 57131 24532 57917 24588
rect 57973 24532 58557 24588
rect 58613 24532 58740 24588
rect 53284 24528 58740 24532
rect 58804 24528 58820 24592
rect 58884 24528 58900 24592
rect 58964 24528 58980 24592
rect 59044 24528 59060 24592
rect 59124 24528 59140 24592
rect 59204 24528 59220 24592
rect 59284 24588 64740 24592
rect 59284 24532 60418 24588
rect 60474 24532 60576 24588
rect 60632 24532 62620 24588
rect 62676 24532 62700 24588
rect 62756 24532 64740 24588
rect 59284 24528 64740 24532
rect 64804 24528 64820 24592
rect 64884 24528 64900 24592
rect 64964 24528 64980 24592
rect 65044 24528 65060 24592
rect 65124 24528 65140 24592
rect 65204 24528 65220 24592
rect 65284 24528 70740 24592
rect 70804 24528 70820 24592
rect 70884 24528 70900 24592
rect 70964 24528 70980 24592
rect 71044 24528 71060 24592
rect 71124 24528 71140 24592
rect 71204 24528 71220 24592
rect 71284 24588 75028 24592
rect 71284 24532 74216 24588
rect 74272 24532 74296 24588
rect 74352 24532 74376 24588
rect 74432 24532 74456 24588
rect 74512 24532 75028 24588
rect 71284 24528 75028 24532
rect 964 24512 75028 24528
rect 964 24508 4740 24512
rect 964 24452 2136 24508
rect 2192 24452 4740 24508
rect 964 24448 4740 24452
rect 4804 24448 4820 24512
rect 4884 24448 4900 24512
rect 4964 24448 4980 24512
rect 5044 24448 5060 24512
rect 5124 24448 5140 24512
rect 5204 24448 5220 24512
rect 5284 24508 10740 24512
rect 5284 24452 5632 24508
rect 5688 24452 8522 24508
rect 8578 24452 10740 24508
rect 5284 24448 10740 24452
rect 10804 24448 10820 24512
rect 10884 24448 10900 24512
rect 10964 24448 10980 24512
rect 11044 24448 11060 24512
rect 11124 24448 11140 24512
rect 11204 24448 11220 24512
rect 11284 24508 16740 24512
rect 11284 24452 11412 24508
rect 11468 24452 14302 24508
rect 14358 24452 16740 24508
rect 11284 24448 16740 24452
rect 16804 24448 16820 24512
rect 16884 24448 16900 24512
rect 16964 24448 16980 24512
rect 17044 24448 17060 24512
rect 17124 24448 17140 24512
rect 17204 24508 17220 24512
rect 17284 24508 22740 24512
rect 17284 24452 20082 24508
rect 20138 24452 22740 24508
rect 17204 24448 17220 24452
rect 17284 24448 22740 24452
rect 22804 24448 22820 24512
rect 22884 24448 22900 24512
rect 22964 24508 22980 24512
rect 22964 24452 22972 24508
rect 22964 24448 22980 24452
rect 23044 24448 23060 24512
rect 23124 24448 23140 24512
rect 23204 24448 23220 24512
rect 23284 24508 28740 24512
rect 28804 24508 28820 24512
rect 23284 24452 25862 24508
rect 25918 24452 28740 24508
rect 28808 24452 28820 24508
rect 23284 24448 28740 24452
rect 28804 24448 28820 24452
rect 28884 24448 28900 24512
rect 28964 24448 28980 24512
rect 29044 24448 29060 24512
rect 29124 24448 29140 24512
rect 29204 24448 29220 24512
rect 29284 24508 34740 24512
rect 29284 24452 31642 24508
rect 31698 24452 34532 24508
rect 34588 24452 34740 24508
rect 29284 24448 34740 24452
rect 34804 24448 34820 24512
rect 34884 24448 34900 24512
rect 34964 24448 34980 24512
rect 35044 24448 35060 24512
rect 35124 24448 35140 24512
rect 35204 24448 35220 24512
rect 35284 24508 40740 24512
rect 35284 24452 37422 24508
rect 37478 24452 40312 24508
rect 40368 24452 40740 24508
rect 35284 24448 40740 24452
rect 40804 24448 40820 24512
rect 40884 24448 40900 24512
rect 40964 24448 40980 24512
rect 41044 24448 41060 24512
rect 41124 24448 41140 24512
rect 41204 24448 41220 24512
rect 41284 24508 46740 24512
rect 41284 24452 43202 24508
rect 43258 24452 46092 24508
rect 46148 24452 46740 24508
rect 41284 24448 46740 24452
rect 46804 24448 46820 24512
rect 46884 24448 46900 24512
rect 46964 24448 46980 24512
rect 47044 24448 47060 24512
rect 47124 24448 47140 24512
rect 47204 24448 47220 24512
rect 47284 24508 52740 24512
rect 47284 24452 49100 24508
rect 49156 24452 52329 24508
rect 52385 24452 52740 24508
rect 47284 24448 52740 24452
rect 52804 24448 52820 24512
rect 52884 24448 52900 24512
rect 52964 24448 52980 24512
rect 53044 24448 53060 24512
rect 53124 24448 53140 24512
rect 53204 24448 53220 24512
rect 53284 24508 58740 24512
rect 53284 24452 53730 24508
rect 53786 24452 53898 24508
rect 53954 24452 54642 24508
rect 54698 24452 55032 24508
rect 55088 24452 55748 24508
rect 55804 24452 56326 24508
rect 56382 24452 56771 24508
rect 56827 24452 57075 24508
rect 57131 24452 57917 24508
rect 57973 24452 58557 24508
rect 58613 24452 58740 24508
rect 53284 24448 58740 24452
rect 58804 24448 58820 24512
rect 58884 24448 58900 24512
rect 58964 24448 58980 24512
rect 59044 24448 59060 24512
rect 59124 24448 59140 24512
rect 59204 24448 59220 24512
rect 59284 24508 64740 24512
rect 59284 24452 60418 24508
rect 60474 24452 60576 24508
rect 60632 24452 62620 24508
rect 62676 24452 62700 24508
rect 62756 24452 64740 24508
rect 59284 24448 64740 24452
rect 64804 24448 64820 24512
rect 64884 24448 64900 24512
rect 64964 24448 64980 24512
rect 65044 24448 65060 24512
rect 65124 24448 65140 24512
rect 65204 24448 65220 24512
rect 65284 24448 70740 24512
rect 70804 24448 70820 24512
rect 70884 24448 70900 24512
rect 70964 24448 70980 24512
rect 71044 24448 71060 24512
rect 71124 24448 71140 24512
rect 71204 24448 71220 24512
rect 71284 24508 75028 24512
rect 71284 24452 74216 24508
rect 74272 24452 74296 24508
rect 74352 24452 74376 24508
rect 74432 24452 74456 24508
rect 74512 24452 75028 24508
rect 71284 24448 75028 24452
rect 964 24432 75028 24448
rect 964 24428 4740 24432
rect 964 24372 2136 24428
rect 2192 24372 4740 24428
rect 964 24368 4740 24372
rect 4804 24368 4820 24432
rect 4884 24368 4900 24432
rect 4964 24368 4980 24432
rect 5044 24368 5060 24432
rect 5124 24368 5140 24432
rect 5204 24368 5220 24432
rect 5284 24428 10740 24432
rect 5284 24372 5632 24428
rect 5688 24372 8522 24428
rect 8578 24372 10740 24428
rect 5284 24368 10740 24372
rect 10804 24368 10820 24432
rect 10884 24368 10900 24432
rect 10964 24368 10980 24432
rect 11044 24368 11060 24432
rect 11124 24368 11140 24432
rect 11204 24368 11220 24432
rect 11284 24428 16740 24432
rect 11284 24372 11412 24428
rect 11468 24372 14302 24428
rect 14358 24372 16740 24428
rect 11284 24368 16740 24372
rect 16804 24368 16820 24432
rect 16884 24368 16900 24432
rect 16964 24368 16980 24432
rect 17044 24368 17060 24432
rect 17124 24368 17140 24432
rect 17204 24428 17220 24432
rect 17284 24428 22740 24432
rect 17284 24372 20082 24428
rect 20138 24372 22740 24428
rect 17204 24368 17220 24372
rect 17284 24368 22740 24372
rect 22804 24368 22820 24432
rect 22884 24368 22900 24432
rect 22964 24428 22980 24432
rect 22964 24372 22972 24428
rect 22964 24368 22980 24372
rect 23044 24368 23060 24432
rect 23124 24368 23140 24432
rect 23204 24368 23220 24432
rect 23284 24428 28740 24432
rect 28804 24428 28820 24432
rect 23284 24372 25862 24428
rect 25918 24372 28740 24428
rect 28808 24372 28820 24428
rect 23284 24368 28740 24372
rect 28804 24368 28820 24372
rect 28884 24368 28900 24432
rect 28964 24368 28980 24432
rect 29044 24368 29060 24432
rect 29124 24368 29140 24432
rect 29204 24368 29220 24432
rect 29284 24428 34740 24432
rect 29284 24372 31642 24428
rect 31698 24372 34532 24428
rect 34588 24372 34740 24428
rect 29284 24368 34740 24372
rect 34804 24368 34820 24432
rect 34884 24368 34900 24432
rect 34964 24368 34980 24432
rect 35044 24368 35060 24432
rect 35124 24368 35140 24432
rect 35204 24368 35220 24432
rect 35284 24428 40740 24432
rect 35284 24372 37422 24428
rect 37478 24372 40312 24428
rect 40368 24372 40740 24428
rect 35284 24368 40740 24372
rect 40804 24368 40820 24432
rect 40884 24368 40900 24432
rect 40964 24368 40980 24432
rect 41044 24368 41060 24432
rect 41124 24368 41140 24432
rect 41204 24368 41220 24432
rect 41284 24428 46740 24432
rect 41284 24372 43202 24428
rect 43258 24372 46092 24428
rect 46148 24372 46740 24428
rect 41284 24368 46740 24372
rect 46804 24368 46820 24432
rect 46884 24368 46900 24432
rect 46964 24368 46980 24432
rect 47044 24368 47060 24432
rect 47124 24368 47140 24432
rect 47204 24368 47220 24432
rect 47284 24428 52740 24432
rect 47284 24372 49100 24428
rect 49156 24372 52329 24428
rect 52385 24372 52740 24428
rect 47284 24368 52740 24372
rect 52804 24368 52820 24432
rect 52884 24368 52900 24432
rect 52964 24368 52980 24432
rect 53044 24368 53060 24432
rect 53124 24368 53140 24432
rect 53204 24368 53220 24432
rect 53284 24428 58740 24432
rect 53284 24372 53730 24428
rect 53786 24372 53898 24428
rect 53954 24372 54642 24428
rect 54698 24372 55032 24428
rect 55088 24372 55748 24428
rect 55804 24372 56326 24428
rect 56382 24372 56771 24428
rect 56827 24372 57075 24428
rect 57131 24372 57917 24428
rect 57973 24372 58557 24428
rect 58613 24372 58740 24428
rect 53284 24368 58740 24372
rect 58804 24368 58820 24432
rect 58884 24368 58900 24432
rect 58964 24368 58980 24432
rect 59044 24368 59060 24432
rect 59124 24368 59140 24432
rect 59204 24368 59220 24432
rect 59284 24428 64740 24432
rect 59284 24372 60418 24428
rect 60474 24372 60576 24428
rect 60632 24372 62620 24428
rect 62676 24372 62700 24428
rect 62756 24372 64740 24428
rect 59284 24368 64740 24372
rect 64804 24368 64820 24432
rect 64884 24368 64900 24432
rect 64964 24368 64980 24432
rect 65044 24368 65060 24432
rect 65124 24368 65140 24432
rect 65204 24368 65220 24432
rect 65284 24368 70740 24432
rect 70804 24368 70820 24432
rect 70884 24368 70900 24432
rect 70964 24368 70980 24432
rect 71044 24368 71060 24432
rect 71124 24368 71140 24432
rect 71204 24368 71220 24432
rect 71284 24428 75028 24432
rect 71284 24372 74216 24428
rect 74272 24372 74296 24428
rect 74352 24372 74376 24428
rect 74432 24372 74456 24428
rect 74512 24372 75028 24428
rect 71284 24368 75028 24372
rect 964 24352 75028 24368
rect 964 24348 4740 24352
rect 964 24292 2136 24348
rect 2192 24292 4740 24348
rect 964 24288 4740 24292
rect 4804 24288 4820 24352
rect 4884 24288 4900 24352
rect 4964 24288 4980 24352
rect 5044 24288 5060 24352
rect 5124 24288 5140 24352
rect 5204 24288 5220 24352
rect 5284 24348 10740 24352
rect 5284 24292 5632 24348
rect 5688 24292 8522 24348
rect 8578 24292 10740 24348
rect 5284 24288 10740 24292
rect 10804 24288 10820 24352
rect 10884 24288 10900 24352
rect 10964 24288 10980 24352
rect 11044 24288 11060 24352
rect 11124 24288 11140 24352
rect 11204 24288 11220 24352
rect 11284 24348 16740 24352
rect 11284 24292 11412 24348
rect 11468 24292 14302 24348
rect 14358 24292 16740 24348
rect 11284 24288 16740 24292
rect 16804 24288 16820 24352
rect 16884 24288 16900 24352
rect 16964 24288 16980 24352
rect 17044 24288 17060 24352
rect 17124 24288 17140 24352
rect 17204 24348 17220 24352
rect 17284 24348 22740 24352
rect 17284 24292 20082 24348
rect 20138 24292 22740 24348
rect 17204 24288 17220 24292
rect 17284 24288 22740 24292
rect 22804 24288 22820 24352
rect 22884 24288 22900 24352
rect 22964 24348 22980 24352
rect 22964 24292 22972 24348
rect 22964 24288 22980 24292
rect 23044 24288 23060 24352
rect 23124 24288 23140 24352
rect 23204 24288 23220 24352
rect 23284 24348 28740 24352
rect 28804 24348 28820 24352
rect 23284 24292 25862 24348
rect 25918 24292 28740 24348
rect 28808 24292 28820 24348
rect 23284 24288 28740 24292
rect 28804 24288 28820 24292
rect 28884 24288 28900 24352
rect 28964 24288 28980 24352
rect 29044 24288 29060 24352
rect 29124 24288 29140 24352
rect 29204 24288 29220 24352
rect 29284 24348 34740 24352
rect 29284 24292 31642 24348
rect 31698 24292 34532 24348
rect 34588 24292 34740 24348
rect 29284 24288 34740 24292
rect 34804 24288 34820 24352
rect 34884 24288 34900 24352
rect 34964 24288 34980 24352
rect 35044 24288 35060 24352
rect 35124 24288 35140 24352
rect 35204 24288 35220 24352
rect 35284 24348 40740 24352
rect 35284 24292 37422 24348
rect 37478 24292 40312 24348
rect 40368 24292 40740 24348
rect 35284 24288 40740 24292
rect 40804 24288 40820 24352
rect 40884 24288 40900 24352
rect 40964 24288 40980 24352
rect 41044 24288 41060 24352
rect 41124 24288 41140 24352
rect 41204 24288 41220 24352
rect 41284 24348 46740 24352
rect 41284 24292 43202 24348
rect 43258 24292 46092 24348
rect 46148 24292 46740 24348
rect 41284 24288 46740 24292
rect 46804 24288 46820 24352
rect 46884 24288 46900 24352
rect 46964 24288 46980 24352
rect 47044 24288 47060 24352
rect 47124 24288 47140 24352
rect 47204 24288 47220 24352
rect 47284 24348 52740 24352
rect 47284 24292 49100 24348
rect 49156 24292 52329 24348
rect 52385 24292 52740 24348
rect 47284 24288 52740 24292
rect 52804 24288 52820 24352
rect 52884 24288 52900 24352
rect 52964 24288 52980 24352
rect 53044 24288 53060 24352
rect 53124 24288 53140 24352
rect 53204 24288 53220 24352
rect 53284 24348 58740 24352
rect 53284 24292 53730 24348
rect 53786 24292 53898 24348
rect 53954 24292 54642 24348
rect 54698 24292 55032 24348
rect 55088 24292 55748 24348
rect 55804 24292 56326 24348
rect 56382 24292 56771 24348
rect 56827 24292 57075 24348
rect 57131 24292 57917 24348
rect 57973 24292 58557 24348
rect 58613 24292 58740 24348
rect 53284 24288 58740 24292
rect 58804 24288 58820 24352
rect 58884 24288 58900 24352
rect 58964 24288 58980 24352
rect 59044 24288 59060 24352
rect 59124 24288 59140 24352
rect 59204 24288 59220 24352
rect 59284 24348 64740 24352
rect 59284 24292 60418 24348
rect 60474 24292 60576 24348
rect 60632 24292 62620 24348
rect 62676 24292 62700 24348
rect 62756 24292 64740 24348
rect 59284 24288 64740 24292
rect 64804 24288 64820 24352
rect 64884 24288 64900 24352
rect 64964 24288 64980 24352
rect 65044 24288 65060 24352
rect 65124 24288 65140 24352
rect 65204 24288 65220 24352
rect 65284 24288 70740 24352
rect 70804 24288 70820 24352
rect 70884 24288 70900 24352
rect 70964 24288 70980 24352
rect 71044 24288 71060 24352
rect 71124 24288 71140 24352
rect 71204 24288 71220 24352
rect 71284 24348 75028 24352
rect 71284 24292 74216 24348
rect 74272 24292 74296 24348
rect 74352 24292 74376 24348
rect 74432 24292 74456 24348
rect 74512 24292 75028 24348
rect 71284 24288 75028 24292
rect 964 24264 75028 24288
rect 67030 23564 67036 23628
rect 67100 23626 67106 23628
rect 67173 23626 67239 23629
rect 67100 23624 67239 23626
rect 67100 23568 67178 23624
rect 67234 23568 67239 23624
rect 67100 23566 67239 23568
rect 67100 23564 67106 23566
rect 67173 23563 67239 23566
rect 67265 23492 67331 23493
rect 67214 23428 67220 23492
rect 67284 23490 67331 23492
rect 67284 23488 67376 23490
rect 67326 23432 67376 23488
rect 67284 23430 67376 23432
rect 67284 23428 67331 23430
rect 67265 23427 67331 23428
rect 66529 22676 66595 22677
rect 66478 22674 66484 22676
rect 66438 22614 66484 22674
rect 66548 22672 66595 22676
rect 66590 22616 66595 22672
rect 66478 22612 66484 22614
rect 66548 22612 66595 22616
rect 66529 22611 66595 22612
rect 66253 22404 66319 22405
rect 66253 22400 66300 22404
rect 66364 22402 66370 22404
rect 66253 22344 66258 22400
rect 66253 22340 66300 22344
rect 66364 22342 66410 22402
rect 66364 22340 66370 22342
rect 66253 22339 66319 22340
rect 964 22240 75028 22264
rect 964 22176 1740 22240
rect 1804 22176 1820 22240
rect 1884 22176 1900 22240
rect 1964 22176 1980 22240
rect 2044 22176 2060 22240
rect 2124 22176 2140 22240
rect 2204 22176 2220 22240
rect 2284 22236 7740 22240
rect 2332 22180 2356 22236
rect 2412 22180 5485 22236
rect 5541 22180 7740 22236
rect 2284 22176 7740 22180
rect 7804 22176 7820 22240
rect 7884 22176 7900 22240
rect 7964 22176 7980 22240
rect 8044 22176 8060 22240
rect 8124 22176 8140 22240
rect 8204 22176 8220 22240
rect 8284 22236 13740 22240
rect 8284 22180 8375 22236
rect 8431 22180 11265 22236
rect 11321 22180 13740 22236
rect 8284 22176 13740 22180
rect 13804 22176 13820 22240
rect 13884 22176 13900 22240
rect 13964 22176 13980 22240
rect 14044 22176 14060 22240
rect 14124 22176 14140 22240
rect 14204 22236 14220 22240
rect 14211 22180 14220 22236
rect 14204 22176 14220 22180
rect 14284 22236 19740 22240
rect 14284 22180 17045 22236
rect 17101 22180 19740 22236
rect 14284 22176 19740 22180
rect 19804 22176 19820 22240
rect 19884 22176 19900 22240
rect 19964 22236 19980 22240
rect 19964 22176 19980 22180
rect 20044 22176 20060 22240
rect 20124 22176 20140 22240
rect 20204 22176 20220 22240
rect 20284 22236 25740 22240
rect 20284 22180 22825 22236
rect 22881 22180 25715 22236
rect 20284 22176 25740 22180
rect 25804 22176 25820 22240
rect 25884 22176 25900 22240
rect 25964 22176 25980 22240
rect 26044 22176 26060 22240
rect 26124 22176 26140 22240
rect 26204 22176 26220 22240
rect 26284 22236 31740 22240
rect 26284 22180 28605 22236
rect 28661 22180 31495 22236
rect 31551 22180 31740 22236
rect 26284 22176 31740 22180
rect 31804 22176 31820 22240
rect 31884 22176 31900 22240
rect 31964 22176 31980 22240
rect 32044 22176 32060 22240
rect 32124 22176 32140 22240
rect 32204 22176 32220 22240
rect 32284 22236 37740 22240
rect 32284 22180 34385 22236
rect 34441 22180 37275 22236
rect 37331 22180 37740 22236
rect 32284 22176 37740 22180
rect 37804 22176 37820 22240
rect 37884 22176 37900 22240
rect 37964 22176 37980 22240
rect 38044 22176 38060 22240
rect 38124 22176 38140 22240
rect 38204 22176 38220 22240
rect 38284 22236 43740 22240
rect 38284 22180 40165 22236
rect 40221 22180 43055 22236
rect 43111 22180 43740 22236
rect 38284 22176 43740 22180
rect 43804 22176 43820 22240
rect 43884 22176 43900 22240
rect 43964 22176 43980 22240
rect 44044 22176 44060 22240
rect 44124 22176 44140 22240
rect 44204 22176 44220 22240
rect 44284 22236 49740 22240
rect 49804 22236 49820 22240
rect 49884 22236 49900 22240
rect 44284 22180 45945 22236
rect 46001 22180 48892 22236
rect 48948 22180 49740 22236
rect 49810 22180 49820 22236
rect 49890 22180 49900 22236
rect 44284 22176 49740 22180
rect 49804 22176 49820 22180
rect 49884 22176 49900 22180
rect 49964 22176 49980 22240
rect 50044 22176 50060 22240
rect 50124 22176 50140 22240
rect 50204 22176 50220 22240
rect 50284 22236 55740 22240
rect 50284 22180 53048 22236
rect 53104 22180 53206 22236
rect 53262 22180 53562 22236
rect 53618 22180 54880 22236
rect 54936 22180 55473 22236
rect 55529 22180 55740 22236
rect 50284 22176 55740 22180
rect 55804 22176 55820 22240
rect 55884 22176 55900 22240
rect 55964 22176 55980 22240
rect 56044 22176 56060 22240
rect 56124 22176 56140 22240
rect 56204 22176 56220 22240
rect 56284 22236 61740 22240
rect 56284 22180 56619 22236
rect 56675 22180 58055 22236
rect 58111 22180 58135 22236
rect 58191 22180 59298 22236
rect 59354 22180 59456 22236
rect 59512 22180 59764 22236
rect 59820 22180 59910 22236
rect 59966 22180 60046 22236
rect 60102 22180 60126 22236
rect 60182 22180 61740 22236
rect 56284 22176 61740 22180
rect 61804 22176 61820 22240
rect 61884 22176 61900 22240
rect 61964 22176 61980 22240
rect 62044 22176 62060 22240
rect 62124 22176 62140 22240
rect 62204 22176 62220 22240
rect 62284 22236 67740 22240
rect 62284 22180 62418 22236
rect 62474 22180 62498 22236
rect 62554 22180 67740 22236
rect 62284 22176 67740 22180
rect 67804 22176 67820 22240
rect 67884 22176 67900 22240
rect 67964 22176 67980 22240
rect 68044 22176 68060 22240
rect 68124 22176 68140 22240
rect 68204 22176 68220 22240
rect 68284 22236 73740 22240
rect 68284 22180 71864 22236
rect 71920 22180 71944 22236
rect 72000 22180 72024 22236
rect 72080 22180 72104 22236
rect 72160 22180 73740 22236
rect 68284 22176 73740 22180
rect 73804 22176 73820 22240
rect 73884 22176 73900 22240
rect 73964 22176 73980 22240
rect 74044 22176 74060 22240
rect 74124 22176 74140 22240
rect 74204 22176 74220 22240
rect 74284 22176 75028 22240
rect 964 22160 75028 22176
rect 964 22096 1740 22160
rect 1804 22096 1820 22160
rect 1884 22096 1900 22160
rect 1964 22096 1980 22160
rect 2044 22096 2060 22160
rect 2124 22096 2140 22160
rect 2204 22096 2220 22160
rect 2284 22156 7740 22160
rect 2332 22100 2356 22156
rect 2412 22100 5485 22156
rect 5541 22100 7740 22156
rect 2284 22096 7740 22100
rect 7804 22096 7820 22160
rect 7884 22096 7900 22160
rect 7964 22096 7980 22160
rect 8044 22096 8060 22160
rect 8124 22096 8140 22160
rect 8204 22096 8220 22160
rect 8284 22156 13740 22160
rect 8284 22100 8375 22156
rect 8431 22100 11265 22156
rect 11321 22100 13740 22156
rect 8284 22096 13740 22100
rect 13804 22096 13820 22160
rect 13884 22096 13900 22160
rect 13964 22096 13980 22160
rect 14044 22096 14060 22160
rect 14124 22096 14140 22160
rect 14204 22156 14220 22160
rect 14211 22100 14220 22156
rect 14204 22096 14220 22100
rect 14284 22156 19740 22160
rect 14284 22100 17045 22156
rect 17101 22100 19740 22156
rect 14284 22096 19740 22100
rect 19804 22096 19820 22160
rect 19884 22096 19900 22160
rect 19964 22156 19980 22160
rect 19964 22096 19980 22100
rect 20044 22096 20060 22160
rect 20124 22096 20140 22160
rect 20204 22096 20220 22160
rect 20284 22156 25740 22160
rect 20284 22100 22825 22156
rect 22881 22100 25715 22156
rect 20284 22096 25740 22100
rect 25804 22096 25820 22160
rect 25884 22096 25900 22160
rect 25964 22096 25980 22160
rect 26044 22096 26060 22160
rect 26124 22096 26140 22160
rect 26204 22096 26220 22160
rect 26284 22156 31740 22160
rect 26284 22100 28605 22156
rect 28661 22100 31495 22156
rect 31551 22100 31740 22156
rect 26284 22096 31740 22100
rect 31804 22096 31820 22160
rect 31884 22096 31900 22160
rect 31964 22096 31980 22160
rect 32044 22096 32060 22160
rect 32124 22096 32140 22160
rect 32204 22096 32220 22160
rect 32284 22156 37740 22160
rect 32284 22100 34385 22156
rect 34441 22100 37275 22156
rect 37331 22100 37740 22156
rect 32284 22096 37740 22100
rect 37804 22096 37820 22160
rect 37884 22096 37900 22160
rect 37964 22096 37980 22160
rect 38044 22096 38060 22160
rect 38124 22096 38140 22160
rect 38204 22096 38220 22160
rect 38284 22156 43740 22160
rect 38284 22100 40165 22156
rect 40221 22100 43055 22156
rect 43111 22100 43740 22156
rect 38284 22096 43740 22100
rect 43804 22096 43820 22160
rect 43884 22096 43900 22160
rect 43964 22096 43980 22160
rect 44044 22096 44060 22160
rect 44124 22096 44140 22160
rect 44204 22096 44220 22160
rect 44284 22156 49740 22160
rect 49804 22156 49820 22160
rect 49884 22156 49900 22160
rect 44284 22100 45945 22156
rect 46001 22100 48892 22156
rect 48948 22100 49740 22156
rect 49810 22100 49820 22156
rect 49890 22100 49900 22156
rect 44284 22096 49740 22100
rect 49804 22096 49820 22100
rect 49884 22096 49900 22100
rect 49964 22096 49980 22160
rect 50044 22096 50060 22160
rect 50124 22096 50140 22160
rect 50204 22096 50220 22160
rect 50284 22156 55740 22160
rect 50284 22100 53048 22156
rect 53104 22100 53206 22156
rect 53262 22100 53562 22156
rect 53618 22100 54880 22156
rect 54936 22100 55473 22156
rect 55529 22100 55740 22156
rect 50284 22096 55740 22100
rect 55804 22096 55820 22160
rect 55884 22096 55900 22160
rect 55964 22096 55980 22160
rect 56044 22096 56060 22160
rect 56124 22096 56140 22160
rect 56204 22096 56220 22160
rect 56284 22156 61740 22160
rect 56284 22100 56619 22156
rect 56675 22100 58055 22156
rect 58111 22100 58135 22156
rect 58191 22100 59298 22156
rect 59354 22100 59456 22156
rect 59512 22100 59764 22156
rect 59820 22100 59910 22156
rect 59966 22100 60046 22156
rect 60102 22100 60126 22156
rect 60182 22100 61740 22156
rect 56284 22096 61740 22100
rect 61804 22096 61820 22160
rect 61884 22096 61900 22160
rect 61964 22096 61980 22160
rect 62044 22096 62060 22160
rect 62124 22096 62140 22160
rect 62204 22096 62220 22160
rect 62284 22156 67740 22160
rect 62284 22100 62418 22156
rect 62474 22100 62498 22156
rect 62554 22100 67740 22156
rect 62284 22096 67740 22100
rect 67804 22096 67820 22160
rect 67884 22096 67900 22160
rect 67964 22096 67980 22160
rect 68044 22096 68060 22160
rect 68124 22096 68140 22160
rect 68204 22096 68220 22160
rect 68284 22156 73740 22160
rect 68284 22100 71864 22156
rect 71920 22100 71944 22156
rect 72000 22100 72024 22156
rect 72080 22100 72104 22156
rect 72160 22100 73740 22156
rect 68284 22096 73740 22100
rect 73804 22096 73820 22160
rect 73884 22096 73900 22160
rect 73964 22096 73980 22160
rect 74044 22096 74060 22160
rect 74124 22096 74140 22160
rect 74204 22096 74220 22160
rect 74284 22096 75028 22160
rect 964 22080 75028 22096
rect 964 22016 1740 22080
rect 1804 22016 1820 22080
rect 1884 22016 1900 22080
rect 1964 22016 1980 22080
rect 2044 22016 2060 22080
rect 2124 22016 2140 22080
rect 2204 22016 2220 22080
rect 2284 22076 7740 22080
rect 2332 22020 2356 22076
rect 2412 22020 5485 22076
rect 5541 22020 7740 22076
rect 2284 22016 7740 22020
rect 7804 22016 7820 22080
rect 7884 22016 7900 22080
rect 7964 22016 7980 22080
rect 8044 22016 8060 22080
rect 8124 22016 8140 22080
rect 8204 22016 8220 22080
rect 8284 22076 13740 22080
rect 8284 22020 8375 22076
rect 8431 22020 11265 22076
rect 11321 22020 13740 22076
rect 8284 22016 13740 22020
rect 13804 22016 13820 22080
rect 13884 22016 13900 22080
rect 13964 22016 13980 22080
rect 14044 22016 14060 22080
rect 14124 22016 14140 22080
rect 14204 22076 14220 22080
rect 14211 22020 14220 22076
rect 14204 22016 14220 22020
rect 14284 22076 19740 22080
rect 14284 22020 17045 22076
rect 17101 22020 19740 22076
rect 14284 22016 19740 22020
rect 19804 22016 19820 22080
rect 19884 22016 19900 22080
rect 19964 22076 19980 22080
rect 19964 22016 19980 22020
rect 20044 22016 20060 22080
rect 20124 22016 20140 22080
rect 20204 22016 20220 22080
rect 20284 22076 25740 22080
rect 20284 22020 22825 22076
rect 22881 22020 25715 22076
rect 20284 22016 25740 22020
rect 25804 22016 25820 22080
rect 25884 22016 25900 22080
rect 25964 22016 25980 22080
rect 26044 22016 26060 22080
rect 26124 22016 26140 22080
rect 26204 22016 26220 22080
rect 26284 22076 31740 22080
rect 26284 22020 28605 22076
rect 28661 22020 31495 22076
rect 31551 22020 31740 22076
rect 26284 22016 31740 22020
rect 31804 22016 31820 22080
rect 31884 22016 31900 22080
rect 31964 22016 31980 22080
rect 32044 22016 32060 22080
rect 32124 22016 32140 22080
rect 32204 22016 32220 22080
rect 32284 22076 37740 22080
rect 32284 22020 34385 22076
rect 34441 22020 37275 22076
rect 37331 22020 37740 22076
rect 32284 22016 37740 22020
rect 37804 22016 37820 22080
rect 37884 22016 37900 22080
rect 37964 22016 37980 22080
rect 38044 22016 38060 22080
rect 38124 22016 38140 22080
rect 38204 22016 38220 22080
rect 38284 22076 43740 22080
rect 38284 22020 40165 22076
rect 40221 22020 43055 22076
rect 43111 22020 43740 22076
rect 38284 22016 43740 22020
rect 43804 22016 43820 22080
rect 43884 22016 43900 22080
rect 43964 22016 43980 22080
rect 44044 22016 44060 22080
rect 44124 22016 44140 22080
rect 44204 22016 44220 22080
rect 44284 22076 49740 22080
rect 49804 22076 49820 22080
rect 49884 22076 49900 22080
rect 44284 22020 45945 22076
rect 46001 22020 48892 22076
rect 48948 22020 49740 22076
rect 49810 22020 49820 22076
rect 49890 22020 49900 22076
rect 44284 22016 49740 22020
rect 49804 22016 49820 22020
rect 49884 22016 49900 22020
rect 49964 22016 49980 22080
rect 50044 22016 50060 22080
rect 50124 22016 50140 22080
rect 50204 22016 50220 22080
rect 50284 22076 55740 22080
rect 50284 22020 53048 22076
rect 53104 22020 53206 22076
rect 53262 22020 53562 22076
rect 53618 22020 54880 22076
rect 54936 22020 55473 22076
rect 55529 22020 55740 22076
rect 50284 22016 55740 22020
rect 55804 22016 55820 22080
rect 55884 22016 55900 22080
rect 55964 22016 55980 22080
rect 56044 22016 56060 22080
rect 56124 22016 56140 22080
rect 56204 22016 56220 22080
rect 56284 22076 61740 22080
rect 56284 22020 56619 22076
rect 56675 22020 58055 22076
rect 58111 22020 58135 22076
rect 58191 22020 59298 22076
rect 59354 22020 59456 22076
rect 59512 22020 59764 22076
rect 59820 22020 59910 22076
rect 59966 22020 60046 22076
rect 60102 22020 60126 22076
rect 60182 22020 61740 22076
rect 56284 22016 61740 22020
rect 61804 22016 61820 22080
rect 61884 22016 61900 22080
rect 61964 22016 61980 22080
rect 62044 22016 62060 22080
rect 62124 22016 62140 22080
rect 62204 22016 62220 22080
rect 62284 22076 67740 22080
rect 62284 22020 62418 22076
rect 62474 22020 62498 22076
rect 62554 22020 67740 22076
rect 62284 22016 67740 22020
rect 67804 22016 67820 22080
rect 67884 22016 67900 22080
rect 67964 22016 67980 22080
rect 68044 22016 68060 22080
rect 68124 22016 68140 22080
rect 68204 22016 68220 22080
rect 68284 22076 73740 22080
rect 68284 22020 71864 22076
rect 71920 22020 71944 22076
rect 72000 22020 72024 22076
rect 72080 22020 72104 22076
rect 72160 22020 73740 22076
rect 68284 22016 73740 22020
rect 73804 22016 73820 22080
rect 73884 22016 73900 22080
rect 73964 22016 73980 22080
rect 74044 22016 74060 22080
rect 74124 22016 74140 22080
rect 74204 22016 74220 22080
rect 74284 22016 75028 22080
rect 964 22000 75028 22016
rect 964 21936 1740 22000
rect 1804 21936 1820 22000
rect 1884 21936 1900 22000
rect 1964 21936 1980 22000
rect 2044 21936 2060 22000
rect 2124 21936 2140 22000
rect 2204 21936 2220 22000
rect 2284 21996 7740 22000
rect 2332 21940 2356 21996
rect 2412 21940 5485 21996
rect 5541 21940 7740 21996
rect 2284 21936 7740 21940
rect 7804 21936 7820 22000
rect 7884 21936 7900 22000
rect 7964 21936 7980 22000
rect 8044 21936 8060 22000
rect 8124 21936 8140 22000
rect 8204 21936 8220 22000
rect 8284 21996 13740 22000
rect 8284 21940 8375 21996
rect 8431 21940 11265 21996
rect 11321 21940 13740 21996
rect 8284 21936 13740 21940
rect 13804 21936 13820 22000
rect 13884 21936 13900 22000
rect 13964 21936 13980 22000
rect 14044 21936 14060 22000
rect 14124 21936 14140 22000
rect 14204 21996 14220 22000
rect 14211 21940 14220 21996
rect 14204 21936 14220 21940
rect 14284 21996 19740 22000
rect 14284 21940 17045 21996
rect 17101 21940 19740 21996
rect 14284 21936 19740 21940
rect 19804 21936 19820 22000
rect 19884 21936 19900 22000
rect 19964 21996 19980 22000
rect 19964 21936 19980 21940
rect 20044 21936 20060 22000
rect 20124 21936 20140 22000
rect 20204 21936 20220 22000
rect 20284 21996 25740 22000
rect 20284 21940 22825 21996
rect 22881 21940 25715 21996
rect 20284 21936 25740 21940
rect 25804 21936 25820 22000
rect 25884 21936 25900 22000
rect 25964 21936 25980 22000
rect 26044 21936 26060 22000
rect 26124 21936 26140 22000
rect 26204 21936 26220 22000
rect 26284 21996 31740 22000
rect 26284 21940 28605 21996
rect 28661 21940 31495 21996
rect 31551 21940 31740 21996
rect 26284 21936 31740 21940
rect 31804 21936 31820 22000
rect 31884 21936 31900 22000
rect 31964 21936 31980 22000
rect 32044 21936 32060 22000
rect 32124 21936 32140 22000
rect 32204 21936 32220 22000
rect 32284 21996 37740 22000
rect 32284 21940 34385 21996
rect 34441 21940 37275 21996
rect 37331 21940 37740 21996
rect 32284 21936 37740 21940
rect 37804 21936 37820 22000
rect 37884 21936 37900 22000
rect 37964 21936 37980 22000
rect 38044 21936 38060 22000
rect 38124 21936 38140 22000
rect 38204 21936 38220 22000
rect 38284 21996 43740 22000
rect 38284 21940 40165 21996
rect 40221 21940 43055 21996
rect 43111 21940 43740 21996
rect 38284 21936 43740 21940
rect 43804 21936 43820 22000
rect 43884 21936 43900 22000
rect 43964 21936 43980 22000
rect 44044 21936 44060 22000
rect 44124 21936 44140 22000
rect 44204 21936 44220 22000
rect 44284 21996 49740 22000
rect 49804 21996 49820 22000
rect 49884 21996 49900 22000
rect 44284 21940 45945 21996
rect 46001 21940 48892 21996
rect 48948 21940 49740 21996
rect 49810 21940 49820 21996
rect 49890 21940 49900 21996
rect 44284 21936 49740 21940
rect 49804 21936 49820 21940
rect 49884 21936 49900 21940
rect 49964 21936 49980 22000
rect 50044 21936 50060 22000
rect 50124 21936 50140 22000
rect 50204 21936 50220 22000
rect 50284 21996 55740 22000
rect 50284 21940 53048 21996
rect 53104 21940 53206 21996
rect 53262 21940 53562 21996
rect 53618 21940 54880 21996
rect 54936 21940 55473 21996
rect 55529 21940 55740 21996
rect 50284 21936 55740 21940
rect 55804 21936 55820 22000
rect 55884 21936 55900 22000
rect 55964 21936 55980 22000
rect 56044 21936 56060 22000
rect 56124 21936 56140 22000
rect 56204 21936 56220 22000
rect 56284 21996 61740 22000
rect 56284 21940 56619 21996
rect 56675 21940 58055 21996
rect 58111 21940 58135 21996
rect 58191 21940 59298 21996
rect 59354 21940 59456 21996
rect 59512 21940 59764 21996
rect 59820 21940 59910 21996
rect 59966 21940 60046 21996
rect 60102 21940 60126 21996
rect 60182 21940 61740 21996
rect 56284 21936 61740 21940
rect 61804 21936 61820 22000
rect 61884 21936 61900 22000
rect 61964 21936 61980 22000
rect 62044 21936 62060 22000
rect 62124 21936 62140 22000
rect 62204 21936 62220 22000
rect 62284 21996 67740 22000
rect 62284 21940 62418 21996
rect 62474 21940 62498 21996
rect 62554 21940 67740 21996
rect 62284 21936 67740 21940
rect 67804 21936 67820 22000
rect 67884 21936 67900 22000
rect 67964 21936 67980 22000
rect 68044 21936 68060 22000
rect 68124 21936 68140 22000
rect 68204 21936 68220 22000
rect 68284 21996 73740 22000
rect 68284 21940 71864 21996
rect 71920 21940 71944 21996
rect 72000 21940 72024 21996
rect 72080 21940 72104 21996
rect 72160 21940 73740 21996
rect 68284 21936 73740 21940
rect 73804 21936 73820 22000
rect 73884 21936 73900 22000
rect 73964 21936 73980 22000
rect 74044 21936 74060 22000
rect 74124 21936 74140 22000
rect 74204 21936 74220 22000
rect 74284 21936 75028 22000
rect 964 21912 75028 21936
rect 63677 18186 63743 18189
rect 64454 18186 64460 18188
rect 63677 18184 64460 18186
rect 63677 18128 63682 18184
rect 63738 18128 64460 18184
rect 63677 18126 64460 18128
rect 63677 18123 63743 18126
rect 64454 18124 64460 18126
rect 64524 18124 64530 18188
rect 63166 15812 63172 15876
rect 63236 15874 63242 15876
rect 63585 15874 63651 15877
rect 63236 15872 63651 15874
rect 63236 15816 63590 15872
rect 63646 15816 63651 15872
rect 63236 15814 63651 15816
rect 63236 15812 63242 15814
rect 63585 15811 63651 15814
rect 964 14592 75028 14616
rect 964 14588 4740 14592
rect 964 14532 2136 14588
rect 2192 14532 4740 14588
rect 964 14528 4740 14532
rect 4804 14528 4820 14592
rect 4884 14528 4900 14592
rect 4964 14528 4980 14592
rect 5044 14528 5060 14592
rect 5124 14528 5140 14592
rect 5204 14528 5220 14592
rect 5284 14588 10740 14592
rect 5284 14532 5632 14588
rect 5688 14532 8522 14588
rect 8578 14532 10740 14588
rect 5284 14528 10740 14532
rect 10804 14528 10820 14592
rect 10884 14528 10900 14592
rect 10964 14528 10980 14592
rect 11044 14528 11060 14592
rect 11124 14528 11140 14592
rect 11204 14528 11220 14592
rect 11284 14588 16740 14592
rect 11284 14532 11412 14588
rect 11468 14532 14302 14588
rect 14358 14532 16740 14588
rect 11284 14528 16740 14532
rect 16804 14528 16820 14592
rect 16884 14528 16900 14592
rect 16964 14528 16980 14592
rect 17044 14528 17060 14592
rect 17124 14528 17140 14592
rect 17204 14588 17220 14592
rect 17284 14588 22740 14592
rect 17284 14532 20082 14588
rect 20138 14532 22740 14588
rect 17204 14528 17220 14532
rect 17284 14528 22740 14532
rect 22804 14528 22820 14592
rect 22884 14528 22900 14592
rect 22964 14588 22980 14592
rect 22964 14532 22972 14588
rect 22964 14528 22980 14532
rect 23044 14528 23060 14592
rect 23124 14528 23140 14592
rect 23204 14528 23220 14592
rect 23284 14588 28740 14592
rect 28804 14588 28820 14592
rect 23284 14532 25862 14588
rect 25918 14532 28740 14588
rect 28808 14532 28820 14588
rect 23284 14528 28740 14532
rect 28804 14528 28820 14532
rect 28884 14528 28900 14592
rect 28964 14528 28980 14592
rect 29044 14528 29060 14592
rect 29124 14528 29140 14592
rect 29204 14528 29220 14592
rect 29284 14588 34740 14592
rect 29284 14532 31642 14588
rect 31698 14532 34532 14588
rect 34588 14532 34740 14588
rect 29284 14528 34740 14532
rect 34804 14528 34820 14592
rect 34884 14528 34900 14592
rect 34964 14528 34980 14592
rect 35044 14528 35060 14592
rect 35124 14528 35140 14592
rect 35204 14528 35220 14592
rect 35284 14588 40740 14592
rect 35284 14532 37422 14588
rect 37478 14532 40312 14588
rect 40368 14532 40740 14588
rect 35284 14528 40740 14532
rect 40804 14528 40820 14592
rect 40884 14528 40900 14592
rect 40964 14528 40980 14592
rect 41044 14528 41060 14592
rect 41124 14528 41140 14592
rect 41204 14528 41220 14592
rect 41284 14588 46740 14592
rect 41284 14532 43202 14588
rect 43258 14532 46092 14588
rect 46148 14532 46740 14588
rect 41284 14528 46740 14532
rect 46804 14528 46820 14592
rect 46884 14528 46900 14592
rect 46964 14528 46980 14592
rect 47044 14528 47060 14592
rect 47124 14528 47140 14592
rect 47204 14528 47220 14592
rect 47284 14588 52740 14592
rect 47284 14532 49100 14588
rect 49156 14532 52329 14588
rect 52385 14532 52740 14588
rect 47284 14528 52740 14532
rect 52804 14528 52820 14592
rect 52884 14528 52900 14592
rect 52964 14528 52980 14592
rect 53044 14528 53060 14592
rect 53124 14528 53140 14592
rect 53204 14528 53220 14592
rect 53284 14588 58740 14592
rect 53284 14532 53730 14588
rect 53786 14532 53898 14588
rect 53954 14532 54642 14588
rect 54698 14532 55032 14588
rect 55088 14532 55748 14588
rect 55804 14532 56326 14588
rect 56382 14532 56771 14588
rect 56827 14532 57075 14588
rect 57131 14532 57917 14588
rect 57973 14532 58557 14588
rect 58613 14532 58740 14588
rect 53284 14528 58740 14532
rect 58804 14528 58820 14592
rect 58884 14528 58900 14592
rect 58964 14528 58980 14592
rect 59044 14528 59060 14592
rect 59124 14528 59140 14592
rect 59204 14528 59220 14592
rect 59284 14588 64740 14592
rect 59284 14532 60418 14588
rect 60474 14532 60576 14588
rect 60632 14532 62620 14588
rect 62676 14532 62700 14588
rect 62756 14532 64740 14588
rect 59284 14528 64740 14532
rect 64804 14528 64820 14592
rect 64884 14528 64900 14592
rect 64964 14528 64980 14592
rect 65044 14528 65060 14592
rect 65124 14528 65140 14592
rect 65204 14528 65220 14592
rect 65284 14528 70740 14592
rect 70804 14528 70820 14592
rect 70884 14528 70900 14592
rect 70964 14528 70980 14592
rect 71044 14528 71060 14592
rect 71124 14528 71140 14592
rect 71204 14528 71220 14592
rect 71284 14588 75028 14592
rect 71284 14532 74216 14588
rect 74272 14532 74296 14588
rect 74352 14532 74376 14588
rect 74432 14532 74456 14588
rect 74512 14532 75028 14588
rect 71284 14528 75028 14532
rect 964 14512 75028 14528
rect 964 14508 4740 14512
rect 964 14452 2136 14508
rect 2192 14452 4740 14508
rect 964 14448 4740 14452
rect 4804 14448 4820 14512
rect 4884 14448 4900 14512
rect 4964 14448 4980 14512
rect 5044 14448 5060 14512
rect 5124 14448 5140 14512
rect 5204 14448 5220 14512
rect 5284 14508 10740 14512
rect 5284 14452 5632 14508
rect 5688 14452 8522 14508
rect 8578 14452 10740 14508
rect 5284 14448 10740 14452
rect 10804 14448 10820 14512
rect 10884 14448 10900 14512
rect 10964 14448 10980 14512
rect 11044 14448 11060 14512
rect 11124 14448 11140 14512
rect 11204 14448 11220 14512
rect 11284 14508 16740 14512
rect 11284 14452 11412 14508
rect 11468 14452 14302 14508
rect 14358 14452 16740 14508
rect 11284 14448 16740 14452
rect 16804 14448 16820 14512
rect 16884 14448 16900 14512
rect 16964 14448 16980 14512
rect 17044 14448 17060 14512
rect 17124 14448 17140 14512
rect 17204 14508 17220 14512
rect 17284 14508 22740 14512
rect 17284 14452 20082 14508
rect 20138 14452 22740 14508
rect 17204 14448 17220 14452
rect 17284 14448 22740 14452
rect 22804 14448 22820 14512
rect 22884 14448 22900 14512
rect 22964 14508 22980 14512
rect 22964 14452 22972 14508
rect 22964 14448 22980 14452
rect 23044 14448 23060 14512
rect 23124 14448 23140 14512
rect 23204 14448 23220 14512
rect 23284 14508 28740 14512
rect 28804 14508 28820 14512
rect 23284 14452 25862 14508
rect 25918 14452 28740 14508
rect 28808 14452 28820 14508
rect 23284 14448 28740 14452
rect 28804 14448 28820 14452
rect 28884 14448 28900 14512
rect 28964 14448 28980 14512
rect 29044 14448 29060 14512
rect 29124 14448 29140 14512
rect 29204 14448 29220 14512
rect 29284 14508 34740 14512
rect 29284 14452 31642 14508
rect 31698 14452 34532 14508
rect 34588 14452 34740 14508
rect 29284 14448 34740 14452
rect 34804 14448 34820 14512
rect 34884 14448 34900 14512
rect 34964 14448 34980 14512
rect 35044 14448 35060 14512
rect 35124 14448 35140 14512
rect 35204 14448 35220 14512
rect 35284 14508 40740 14512
rect 35284 14452 37422 14508
rect 37478 14452 40312 14508
rect 40368 14452 40740 14508
rect 35284 14448 40740 14452
rect 40804 14448 40820 14512
rect 40884 14448 40900 14512
rect 40964 14448 40980 14512
rect 41044 14448 41060 14512
rect 41124 14448 41140 14512
rect 41204 14448 41220 14512
rect 41284 14508 46740 14512
rect 41284 14452 43202 14508
rect 43258 14452 46092 14508
rect 46148 14452 46740 14508
rect 41284 14448 46740 14452
rect 46804 14448 46820 14512
rect 46884 14448 46900 14512
rect 46964 14448 46980 14512
rect 47044 14448 47060 14512
rect 47124 14448 47140 14512
rect 47204 14448 47220 14512
rect 47284 14508 52740 14512
rect 47284 14452 49100 14508
rect 49156 14452 52329 14508
rect 52385 14452 52740 14508
rect 47284 14448 52740 14452
rect 52804 14448 52820 14512
rect 52884 14448 52900 14512
rect 52964 14448 52980 14512
rect 53044 14448 53060 14512
rect 53124 14448 53140 14512
rect 53204 14448 53220 14512
rect 53284 14508 58740 14512
rect 53284 14452 53730 14508
rect 53786 14452 53898 14508
rect 53954 14452 54642 14508
rect 54698 14452 55032 14508
rect 55088 14452 55748 14508
rect 55804 14452 56326 14508
rect 56382 14452 56771 14508
rect 56827 14452 57075 14508
rect 57131 14452 57917 14508
rect 57973 14452 58557 14508
rect 58613 14452 58740 14508
rect 53284 14448 58740 14452
rect 58804 14448 58820 14512
rect 58884 14448 58900 14512
rect 58964 14448 58980 14512
rect 59044 14448 59060 14512
rect 59124 14448 59140 14512
rect 59204 14448 59220 14512
rect 59284 14508 64740 14512
rect 59284 14452 60418 14508
rect 60474 14452 60576 14508
rect 60632 14452 62620 14508
rect 62676 14452 62700 14508
rect 62756 14452 64740 14508
rect 59284 14448 64740 14452
rect 64804 14448 64820 14512
rect 64884 14448 64900 14512
rect 64964 14448 64980 14512
rect 65044 14448 65060 14512
rect 65124 14448 65140 14512
rect 65204 14448 65220 14512
rect 65284 14448 70740 14512
rect 70804 14448 70820 14512
rect 70884 14448 70900 14512
rect 70964 14448 70980 14512
rect 71044 14448 71060 14512
rect 71124 14448 71140 14512
rect 71204 14448 71220 14512
rect 71284 14508 75028 14512
rect 71284 14452 74216 14508
rect 74272 14452 74296 14508
rect 74352 14452 74376 14508
rect 74432 14452 74456 14508
rect 74512 14452 75028 14508
rect 71284 14448 75028 14452
rect 964 14432 75028 14448
rect 964 14428 4740 14432
rect 964 14372 2136 14428
rect 2192 14372 4740 14428
rect 964 14368 4740 14372
rect 4804 14368 4820 14432
rect 4884 14368 4900 14432
rect 4964 14368 4980 14432
rect 5044 14368 5060 14432
rect 5124 14368 5140 14432
rect 5204 14368 5220 14432
rect 5284 14428 10740 14432
rect 5284 14372 5632 14428
rect 5688 14372 8522 14428
rect 8578 14372 10740 14428
rect 5284 14368 10740 14372
rect 10804 14368 10820 14432
rect 10884 14368 10900 14432
rect 10964 14368 10980 14432
rect 11044 14368 11060 14432
rect 11124 14368 11140 14432
rect 11204 14368 11220 14432
rect 11284 14428 16740 14432
rect 11284 14372 11412 14428
rect 11468 14372 14302 14428
rect 14358 14372 16740 14428
rect 11284 14368 16740 14372
rect 16804 14368 16820 14432
rect 16884 14368 16900 14432
rect 16964 14368 16980 14432
rect 17044 14368 17060 14432
rect 17124 14368 17140 14432
rect 17204 14428 17220 14432
rect 17284 14428 22740 14432
rect 17284 14372 20082 14428
rect 20138 14372 22740 14428
rect 17204 14368 17220 14372
rect 17284 14368 22740 14372
rect 22804 14368 22820 14432
rect 22884 14368 22900 14432
rect 22964 14428 22980 14432
rect 22964 14372 22972 14428
rect 22964 14368 22980 14372
rect 23044 14368 23060 14432
rect 23124 14368 23140 14432
rect 23204 14368 23220 14432
rect 23284 14428 28740 14432
rect 28804 14428 28820 14432
rect 23284 14372 25862 14428
rect 25918 14372 28740 14428
rect 28808 14372 28820 14428
rect 23284 14368 28740 14372
rect 28804 14368 28820 14372
rect 28884 14368 28900 14432
rect 28964 14368 28980 14432
rect 29044 14368 29060 14432
rect 29124 14368 29140 14432
rect 29204 14368 29220 14432
rect 29284 14428 34740 14432
rect 29284 14372 31642 14428
rect 31698 14372 34532 14428
rect 34588 14372 34740 14428
rect 29284 14368 34740 14372
rect 34804 14368 34820 14432
rect 34884 14368 34900 14432
rect 34964 14368 34980 14432
rect 35044 14368 35060 14432
rect 35124 14368 35140 14432
rect 35204 14368 35220 14432
rect 35284 14428 40740 14432
rect 35284 14372 37422 14428
rect 37478 14372 40312 14428
rect 40368 14372 40740 14428
rect 35284 14368 40740 14372
rect 40804 14368 40820 14432
rect 40884 14368 40900 14432
rect 40964 14368 40980 14432
rect 41044 14368 41060 14432
rect 41124 14368 41140 14432
rect 41204 14368 41220 14432
rect 41284 14428 46740 14432
rect 41284 14372 43202 14428
rect 43258 14372 46092 14428
rect 46148 14372 46740 14428
rect 41284 14368 46740 14372
rect 46804 14368 46820 14432
rect 46884 14368 46900 14432
rect 46964 14368 46980 14432
rect 47044 14368 47060 14432
rect 47124 14368 47140 14432
rect 47204 14368 47220 14432
rect 47284 14428 52740 14432
rect 47284 14372 49100 14428
rect 49156 14372 52329 14428
rect 52385 14372 52740 14428
rect 47284 14368 52740 14372
rect 52804 14368 52820 14432
rect 52884 14368 52900 14432
rect 52964 14368 52980 14432
rect 53044 14368 53060 14432
rect 53124 14368 53140 14432
rect 53204 14368 53220 14432
rect 53284 14428 58740 14432
rect 53284 14372 53730 14428
rect 53786 14372 53898 14428
rect 53954 14372 54642 14428
rect 54698 14372 55032 14428
rect 55088 14372 55748 14428
rect 55804 14372 56326 14428
rect 56382 14372 56771 14428
rect 56827 14372 57075 14428
rect 57131 14372 57917 14428
rect 57973 14372 58557 14428
rect 58613 14372 58740 14428
rect 53284 14368 58740 14372
rect 58804 14368 58820 14432
rect 58884 14368 58900 14432
rect 58964 14368 58980 14432
rect 59044 14368 59060 14432
rect 59124 14368 59140 14432
rect 59204 14368 59220 14432
rect 59284 14428 64740 14432
rect 59284 14372 60418 14428
rect 60474 14372 60576 14428
rect 60632 14372 62620 14428
rect 62676 14372 62700 14428
rect 62756 14372 64740 14428
rect 59284 14368 64740 14372
rect 64804 14368 64820 14432
rect 64884 14368 64900 14432
rect 64964 14368 64980 14432
rect 65044 14368 65060 14432
rect 65124 14368 65140 14432
rect 65204 14368 65220 14432
rect 65284 14368 70740 14432
rect 70804 14368 70820 14432
rect 70884 14368 70900 14432
rect 70964 14368 70980 14432
rect 71044 14368 71060 14432
rect 71124 14368 71140 14432
rect 71204 14368 71220 14432
rect 71284 14428 75028 14432
rect 71284 14372 74216 14428
rect 74272 14372 74296 14428
rect 74352 14372 74376 14428
rect 74432 14372 74456 14428
rect 74512 14372 75028 14428
rect 71284 14368 75028 14372
rect 964 14352 75028 14368
rect 964 14348 4740 14352
rect 964 14292 2136 14348
rect 2192 14292 4740 14348
rect 964 14288 4740 14292
rect 4804 14288 4820 14352
rect 4884 14288 4900 14352
rect 4964 14288 4980 14352
rect 5044 14288 5060 14352
rect 5124 14288 5140 14352
rect 5204 14288 5220 14352
rect 5284 14348 10740 14352
rect 5284 14292 5632 14348
rect 5688 14292 8522 14348
rect 8578 14292 10740 14348
rect 5284 14288 10740 14292
rect 10804 14288 10820 14352
rect 10884 14288 10900 14352
rect 10964 14288 10980 14352
rect 11044 14288 11060 14352
rect 11124 14288 11140 14352
rect 11204 14288 11220 14352
rect 11284 14348 16740 14352
rect 11284 14292 11412 14348
rect 11468 14292 14302 14348
rect 14358 14292 16740 14348
rect 11284 14288 16740 14292
rect 16804 14288 16820 14352
rect 16884 14288 16900 14352
rect 16964 14288 16980 14352
rect 17044 14288 17060 14352
rect 17124 14288 17140 14352
rect 17204 14348 17220 14352
rect 17284 14348 22740 14352
rect 17284 14292 20082 14348
rect 20138 14292 22740 14348
rect 17204 14288 17220 14292
rect 17284 14288 22740 14292
rect 22804 14288 22820 14352
rect 22884 14288 22900 14352
rect 22964 14348 22980 14352
rect 22964 14292 22972 14348
rect 22964 14288 22980 14292
rect 23044 14288 23060 14352
rect 23124 14288 23140 14352
rect 23204 14288 23220 14352
rect 23284 14348 28740 14352
rect 28804 14348 28820 14352
rect 23284 14292 25862 14348
rect 25918 14292 28740 14348
rect 28808 14292 28820 14348
rect 23284 14288 28740 14292
rect 28804 14288 28820 14292
rect 28884 14288 28900 14352
rect 28964 14288 28980 14352
rect 29044 14288 29060 14352
rect 29124 14288 29140 14352
rect 29204 14288 29220 14352
rect 29284 14348 34740 14352
rect 29284 14292 31642 14348
rect 31698 14292 34532 14348
rect 34588 14292 34740 14348
rect 29284 14288 34740 14292
rect 34804 14288 34820 14352
rect 34884 14288 34900 14352
rect 34964 14288 34980 14352
rect 35044 14288 35060 14352
rect 35124 14288 35140 14352
rect 35204 14288 35220 14352
rect 35284 14348 40740 14352
rect 35284 14292 37422 14348
rect 37478 14292 40312 14348
rect 40368 14292 40740 14348
rect 35284 14288 40740 14292
rect 40804 14288 40820 14352
rect 40884 14288 40900 14352
rect 40964 14288 40980 14352
rect 41044 14288 41060 14352
rect 41124 14288 41140 14352
rect 41204 14288 41220 14352
rect 41284 14348 46740 14352
rect 41284 14292 43202 14348
rect 43258 14292 46092 14348
rect 46148 14292 46740 14348
rect 41284 14288 46740 14292
rect 46804 14288 46820 14352
rect 46884 14288 46900 14352
rect 46964 14288 46980 14352
rect 47044 14288 47060 14352
rect 47124 14288 47140 14352
rect 47204 14288 47220 14352
rect 47284 14348 52740 14352
rect 47284 14292 49100 14348
rect 49156 14292 52329 14348
rect 52385 14292 52740 14348
rect 47284 14288 52740 14292
rect 52804 14288 52820 14352
rect 52884 14288 52900 14352
rect 52964 14288 52980 14352
rect 53044 14288 53060 14352
rect 53124 14288 53140 14352
rect 53204 14288 53220 14352
rect 53284 14348 58740 14352
rect 53284 14292 53730 14348
rect 53786 14292 53898 14348
rect 53954 14292 54642 14348
rect 54698 14292 55032 14348
rect 55088 14292 55748 14348
rect 55804 14292 56326 14348
rect 56382 14292 56771 14348
rect 56827 14292 57075 14348
rect 57131 14292 57917 14348
rect 57973 14292 58557 14348
rect 58613 14292 58740 14348
rect 53284 14288 58740 14292
rect 58804 14288 58820 14352
rect 58884 14288 58900 14352
rect 58964 14288 58980 14352
rect 59044 14288 59060 14352
rect 59124 14288 59140 14352
rect 59204 14288 59220 14352
rect 59284 14348 64740 14352
rect 59284 14292 60418 14348
rect 60474 14292 60576 14348
rect 60632 14292 62620 14348
rect 62676 14292 62700 14348
rect 62756 14292 64740 14348
rect 59284 14288 64740 14292
rect 64804 14288 64820 14352
rect 64884 14288 64900 14352
rect 64964 14288 64980 14352
rect 65044 14288 65060 14352
rect 65124 14288 65140 14352
rect 65204 14288 65220 14352
rect 65284 14288 70740 14352
rect 70804 14288 70820 14352
rect 70884 14288 70900 14352
rect 70964 14288 70980 14352
rect 71044 14288 71060 14352
rect 71124 14288 71140 14352
rect 71204 14288 71220 14352
rect 71284 14348 75028 14352
rect 71284 14292 74216 14348
rect 74272 14292 74296 14348
rect 74352 14292 74376 14348
rect 74432 14292 74456 14348
rect 74512 14292 75028 14348
rect 71284 14288 75028 14292
rect 964 14264 75028 14288
rect 65926 12684 65932 12748
rect 65996 12746 66002 12748
rect 66069 12746 66135 12749
rect 65996 12744 66135 12746
rect 65996 12688 66074 12744
rect 66130 12688 66135 12744
rect 65996 12686 66135 12688
rect 65996 12684 66002 12686
rect 66069 12683 66135 12686
rect 964 12240 75028 12264
rect 964 12176 1740 12240
rect 1804 12176 1820 12240
rect 1884 12176 1900 12240
rect 1964 12176 1980 12240
rect 2044 12176 2060 12240
rect 2124 12176 2140 12240
rect 2204 12176 2220 12240
rect 2284 12236 7740 12240
rect 2332 12180 2356 12236
rect 2412 12180 5485 12236
rect 5541 12180 7740 12236
rect 2284 12176 7740 12180
rect 7804 12176 7820 12240
rect 7884 12176 7900 12240
rect 7964 12176 7980 12240
rect 8044 12176 8060 12240
rect 8124 12176 8140 12240
rect 8204 12176 8220 12240
rect 8284 12236 13740 12240
rect 8284 12180 8375 12236
rect 8431 12180 11265 12236
rect 11321 12180 13740 12236
rect 8284 12176 13740 12180
rect 13804 12176 13820 12240
rect 13884 12176 13900 12240
rect 13964 12176 13980 12240
rect 14044 12176 14060 12240
rect 14124 12176 14140 12240
rect 14204 12236 14220 12240
rect 14211 12180 14220 12236
rect 14204 12176 14220 12180
rect 14284 12236 19740 12240
rect 14284 12180 17045 12236
rect 17101 12180 19740 12236
rect 14284 12176 19740 12180
rect 19804 12176 19820 12240
rect 19884 12176 19900 12240
rect 19964 12236 19980 12240
rect 19964 12176 19980 12180
rect 20044 12176 20060 12240
rect 20124 12176 20140 12240
rect 20204 12176 20220 12240
rect 20284 12236 25740 12240
rect 20284 12180 22825 12236
rect 22881 12180 25715 12236
rect 20284 12176 25740 12180
rect 25804 12176 25820 12240
rect 25884 12176 25900 12240
rect 25964 12176 25980 12240
rect 26044 12176 26060 12240
rect 26124 12176 26140 12240
rect 26204 12176 26220 12240
rect 26284 12236 31740 12240
rect 26284 12180 28605 12236
rect 28661 12180 31495 12236
rect 31551 12180 31740 12236
rect 26284 12176 31740 12180
rect 31804 12176 31820 12240
rect 31884 12176 31900 12240
rect 31964 12176 31980 12240
rect 32044 12176 32060 12240
rect 32124 12176 32140 12240
rect 32204 12176 32220 12240
rect 32284 12236 37740 12240
rect 32284 12180 34385 12236
rect 34441 12180 37275 12236
rect 37331 12180 37740 12236
rect 32284 12176 37740 12180
rect 37804 12176 37820 12240
rect 37884 12176 37900 12240
rect 37964 12176 37980 12240
rect 38044 12176 38060 12240
rect 38124 12176 38140 12240
rect 38204 12176 38220 12240
rect 38284 12236 43740 12240
rect 38284 12180 40165 12236
rect 40221 12180 43055 12236
rect 43111 12180 43740 12236
rect 38284 12176 43740 12180
rect 43804 12176 43820 12240
rect 43884 12176 43900 12240
rect 43964 12176 43980 12240
rect 44044 12176 44060 12240
rect 44124 12176 44140 12240
rect 44204 12176 44220 12240
rect 44284 12236 49740 12240
rect 49804 12236 49820 12240
rect 49884 12236 49900 12240
rect 44284 12180 45945 12236
rect 46001 12180 48892 12236
rect 48948 12180 49740 12236
rect 49810 12180 49820 12236
rect 49890 12180 49900 12236
rect 44284 12176 49740 12180
rect 49804 12176 49820 12180
rect 49884 12176 49900 12180
rect 49964 12176 49980 12240
rect 50044 12176 50060 12240
rect 50124 12176 50140 12240
rect 50204 12176 50220 12240
rect 50284 12236 55740 12240
rect 50284 12180 53048 12236
rect 53104 12180 53206 12236
rect 53262 12180 53562 12236
rect 53618 12180 54880 12236
rect 54936 12180 55473 12236
rect 55529 12180 55740 12236
rect 50284 12176 55740 12180
rect 55804 12176 55820 12240
rect 55884 12176 55900 12240
rect 55964 12176 55980 12240
rect 56044 12176 56060 12240
rect 56124 12176 56140 12240
rect 56204 12176 56220 12240
rect 56284 12236 61740 12240
rect 56284 12180 56619 12236
rect 56675 12180 58055 12236
rect 58111 12180 58135 12236
rect 58191 12180 59298 12236
rect 59354 12180 59456 12236
rect 59512 12180 59764 12236
rect 59820 12180 59910 12236
rect 59966 12180 60046 12236
rect 60102 12180 60126 12236
rect 60182 12180 61740 12236
rect 56284 12176 61740 12180
rect 61804 12176 61820 12240
rect 61884 12176 61900 12240
rect 61964 12176 61980 12240
rect 62044 12176 62060 12240
rect 62124 12176 62140 12240
rect 62204 12176 62220 12240
rect 62284 12236 67740 12240
rect 62284 12180 62418 12236
rect 62474 12180 62498 12236
rect 62554 12180 67740 12236
rect 62284 12176 67740 12180
rect 67804 12176 67820 12240
rect 67884 12176 67900 12240
rect 67964 12176 67980 12240
rect 68044 12176 68060 12240
rect 68124 12176 68140 12240
rect 68204 12176 68220 12240
rect 68284 12236 73740 12240
rect 68284 12180 71864 12236
rect 71920 12180 71944 12236
rect 72000 12180 72024 12236
rect 72080 12180 72104 12236
rect 72160 12180 73740 12236
rect 68284 12176 73740 12180
rect 73804 12176 73820 12240
rect 73884 12176 73900 12240
rect 73964 12176 73980 12240
rect 74044 12176 74060 12240
rect 74124 12176 74140 12240
rect 74204 12176 74220 12240
rect 74284 12176 75028 12240
rect 964 12160 75028 12176
rect 964 12096 1740 12160
rect 1804 12096 1820 12160
rect 1884 12096 1900 12160
rect 1964 12096 1980 12160
rect 2044 12096 2060 12160
rect 2124 12096 2140 12160
rect 2204 12096 2220 12160
rect 2284 12156 7740 12160
rect 2332 12100 2356 12156
rect 2412 12100 5485 12156
rect 5541 12100 7740 12156
rect 2284 12096 7740 12100
rect 7804 12096 7820 12160
rect 7884 12096 7900 12160
rect 7964 12096 7980 12160
rect 8044 12096 8060 12160
rect 8124 12096 8140 12160
rect 8204 12096 8220 12160
rect 8284 12156 13740 12160
rect 8284 12100 8375 12156
rect 8431 12100 11265 12156
rect 11321 12100 13740 12156
rect 8284 12096 13740 12100
rect 13804 12096 13820 12160
rect 13884 12096 13900 12160
rect 13964 12096 13980 12160
rect 14044 12096 14060 12160
rect 14124 12096 14140 12160
rect 14204 12156 14220 12160
rect 14211 12100 14220 12156
rect 14204 12096 14220 12100
rect 14284 12156 19740 12160
rect 14284 12100 17045 12156
rect 17101 12100 19740 12156
rect 14284 12096 19740 12100
rect 19804 12096 19820 12160
rect 19884 12096 19900 12160
rect 19964 12156 19980 12160
rect 19964 12096 19980 12100
rect 20044 12096 20060 12160
rect 20124 12096 20140 12160
rect 20204 12096 20220 12160
rect 20284 12156 25740 12160
rect 20284 12100 22825 12156
rect 22881 12100 25715 12156
rect 20284 12096 25740 12100
rect 25804 12096 25820 12160
rect 25884 12096 25900 12160
rect 25964 12096 25980 12160
rect 26044 12096 26060 12160
rect 26124 12096 26140 12160
rect 26204 12096 26220 12160
rect 26284 12156 31740 12160
rect 26284 12100 28605 12156
rect 28661 12100 31495 12156
rect 31551 12100 31740 12156
rect 26284 12096 31740 12100
rect 31804 12096 31820 12160
rect 31884 12096 31900 12160
rect 31964 12096 31980 12160
rect 32044 12096 32060 12160
rect 32124 12096 32140 12160
rect 32204 12096 32220 12160
rect 32284 12156 37740 12160
rect 32284 12100 34385 12156
rect 34441 12100 37275 12156
rect 37331 12100 37740 12156
rect 32284 12096 37740 12100
rect 37804 12096 37820 12160
rect 37884 12096 37900 12160
rect 37964 12096 37980 12160
rect 38044 12096 38060 12160
rect 38124 12096 38140 12160
rect 38204 12096 38220 12160
rect 38284 12156 43740 12160
rect 38284 12100 40165 12156
rect 40221 12100 43055 12156
rect 43111 12100 43740 12156
rect 38284 12096 43740 12100
rect 43804 12096 43820 12160
rect 43884 12096 43900 12160
rect 43964 12096 43980 12160
rect 44044 12096 44060 12160
rect 44124 12096 44140 12160
rect 44204 12096 44220 12160
rect 44284 12156 49740 12160
rect 49804 12156 49820 12160
rect 49884 12156 49900 12160
rect 44284 12100 45945 12156
rect 46001 12100 48892 12156
rect 48948 12100 49740 12156
rect 49810 12100 49820 12156
rect 49890 12100 49900 12156
rect 44284 12096 49740 12100
rect 49804 12096 49820 12100
rect 49884 12096 49900 12100
rect 49964 12096 49980 12160
rect 50044 12096 50060 12160
rect 50124 12096 50140 12160
rect 50204 12096 50220 12160
rect 50284 12156 55740 12160
rect 50284 12100 53048 12156
rect 53104 12100 53206 12156
rect 53262 12100 53562 12156
rect 53618 12100 54880 12156
rect 54936 12100 55473 12156
rect 55529 12100 55740 12156
rect 50284 12096 55740 12100
rect 55804 12096 55820 12160
rect 55884 12096 55900 12160
rect 55964 12096 55980 12160
rect 56044 12096 56060 12160
rect 56124 12096 56140 12160
rect 56204 12096 56220 12160
rect 56284 12156 61740 12160
rect 56284 12100 56619 12156
rect 56675 12100 58055 12156
rect 58111 12100 58135 12156
rect 58191 12100 59298 12156
rect 59354 12100 59456 12156
rect 59512 12100 59764 12156
rect 59820 12100 59910 12156
rect 59966 12100 60046 12156
rect 60102 12100 60126 12156
rect 60182 12100 61740 12156
rect 56284 12096 61740 12100
rect 61804 12096 61820 12160
rect 61884 12096 61900 12160
rect 61964 12096 61980 12160
rect 62044 12096 62060 12160
rect 62124 12096 62140 12160
rect 62204 12096 62220 12160
rect 62284 12156 67740 12160
rect 62284 12100 62418 12156
rect 62474 12100 62498 12156
rect 62554 12100 67740 12156
rect 62284 12096 67740 12100
rect 67804 12096 67820 12160
rect 67884 12096 67900 12160
rect 67964 12096 67980 12160
rect 68044 12096 68060 12160
rect 68124 12096 68140 12160
rect 68204 12096 68220 12160
rect 68284 12156 73740 12160
rect 68284 12100 71864 12156
rect 71920 12100 71944 12156
rect 72000 12100 72024 12156
rect 72080 12100 72104 12156
rect 72160 12100 73740 12156
rect 68284 12096 73740 12100
rect 73804 12096 73820 12160
rect 73884 12096 73900 12160
rect 73964 12096 73980 12160
rect 74044 12096 74060 12160
rect 74124 12096 74140 12160
rect 74204 12096 74220 12160
rect 74284 12096 75028 12160
rect 964 12080 75028 12096
rect 964 12016 1740 12080
rect 1804 12016 1820 12080
rect 1884 12016 1900 12080
rect 1964 12016 1980 12080
rect 2044 12016 2060 12080
rect 2124 12016 2140 12080
rect 2204 12016 2220 12080
rect 2284 12076 7740 12080
rect 2332 12020 2356 12076
rect 2412 12020 5485 12076
rect 5541 12020 7740 12076
rect 2284 12016 7740 12020
rect 7804 12016 7820 12080
rect 7884 12016 7900 12080
rect 7964 12016 7980 12080
rect 8044 12016 8060 12080
rect 8124 12016 8140 12080
rect 8204 12016 8220 12080
rect 8284 12076 13740 12080
rect 8284 12020 8375 12076
rect 8431 12020 11265 12076
rect 11321 12020 13740 12076
rect 8284 12016 13740 12020
rect 13804 12016 13820 12080
rect 13884 12016 13900 12080
rect 13964 12016 13980 12080
rect 14044 12016 14060 12080
rect 14124 12016 14140 12080
rect 14204 12076 14220 12080
rect 14211 12020 14220 12076
rect 14204 12016 14220 12020
rect 14284 12076 19740 12080
rect 14284 12020 17045 12076
rect 17101 12020 19740 12076
rect 14284 12016 19740 12020
rect 19804 12016 19820 12080
rect 19884 12016 19900 12080
rect 19964 12076 19980 12080
rect 19964 12016 19980 12020
rect 20044 12016 20060 12080
rect 20124 12016 20140 12080
rect 20204 12016 20220 12080
rect 20284 12076 25740 12080
rect 20284 12020 22825 12076
rect 22881 12020 25715 12076
rect 20284 12016 25740 12020
rect 25804 12016 25820 12080
rect 25884 12016 25900 12080
rect 25964 12016 25980 12080
rect 26044 12016 26060 12080
rect 26124 12016 26140 12080
rect 26204 12016 26220 12080
rect 26284 12076 31740 12080
rect 26284 12020 28605 12076
rect 28661 12020 31495 12076
rect 31551 12020 31740 12076
rect 26284 12016 31740 12020
rect 31804 12016 31820 12080
rect 31884 12016 31900 12080
rect 31964 12016 31980 12080
rect 32044 12016 32060 12080
rect 32124 12016 32140 12080
rect 32204 12016 32220 12080
rect 32284 12076 37740 12080
rect 32284 12020 34385 12076
rect 34441 12020 37275 12076
rect 37331 12020 37740 12076
rect 32284 12016 37740 12020
rect 37804 12016 37820 12080
rect 37884 12016 37900 12080
rect 37964 12016 37980 12080
rect 38044 12016 38060 12080
rect 38124 12016 38140 12080
rect 38204 12016 38220 12080
rect 38284 12076 43740 12080
rect 38284 12020 40165 12076
rect 40221 12020 43055 12076
rect 43111 12020 43740 12076
rect 38284 12016 43740 12020
rect 43804 12016 43820 12080
rect 43884 12016 43900 12080
rect 43964 12016 43980 12080
rect 44044 12016 44060 12080
rect 44124 12016 44140 12080
rect 44204 12016 44220 12080
rect 44284 12076 49740 12080
rect 49804 12076 49820 12080
rect 49884 12076 49900 12080
rect 44284 12020 45945 12076
rect 46001 12020 48892 12076
rect 48948 12020 49740 12076
rect 49810 12020 49820 12076
rect 49890 12020 49900 12076
rect 44284 12016 49740 12020
rect 49804 12016 49820 12020
rect 49884 12016 49900 12020
rect 49964 12016 49980 12080
rect 50044 12016 50060 12080
rect 50124 12016 50140 12080
rect 50204 12016 50220 12080
rect 50284 12076 55740 12080
rect 50284 12020 53048 12076
rect 53104 12020 53206 12076
rect 53262 12020 53562 12076
rect 53618 12020 54880 12076
rect 54936 12020 55473 12076
rect 55529 12020 55740 12076
rect 50284 12016 55740 12020
rect 55804 12016 55820 12080
rect 55884 12016 55900 12080
rect 55964 12016 55980 12080
rect 56044 12016 56060 12080
rect 56124 12016 56140 12080
rect 56204 12016 56220 12080
rect 56284 12076 61740 12080
rect 56284 12020 56619 12076
rect 56675 12020 58055 12076
rect 58111 12020 58135 12076
rect 58191 12020 59298 12076
rect 59354 12020 59456 12076
rect 59512 12020 59764 12076
rect 59820 12020 59910 12076
rect 59966 12020 60046 12076
rect 60102 12020 60126 12076
rect 60182 12020 61740 12076
rect 56284 12016 61740 12020
rect 61804 12016 61820 12080
rect 61884 12016 61900 12080
rect 61964 12016 61980 12080
rect 62044 12016 62060 12080
rect 62124 12016 62140 12080
rect 62204 12016 62220 12080
rect 62284 12076 67740 12080
rect 62284 12020 62418 12076
rect 62474 12020 62498 12076
rect 62554 12020 67740 12076
rect 62284 12016 67740 12020
rect 67804 12016 67820 12080
rect 67884 12016 67900 12080
rect 67964 12016 67980 12080
rect 68044 12016 68060 12080
rect 68124 12016 68140 12080
rect 68204 12016 68220 12080
rect 68284 12076 73740 12080
rect 68284 12020 71864 12076
rect 71920 12020 71944 12076
rect 72000 12020 72024 12076
rect 72080 12020 72104 12076
rect 72160 12020 73740 12076
rect 68284 12016 73740 12020
rect 73804 12016 73820 12080
rect 73884 12016 73900 12080
rect 73964 12016 73980 12080
rect 74044 12016 74060 12080
rect 74124 12016 74140 12080
rect 74204 12016 74220 12080
rect 74284 12016 75028 12080
rect 964 12000 75028 12016
rect 964 11936 1740 12000
rect 1804 11936 1820 12000
rect 1884 11936 1900 12000
rect 1964 11936 1980 12000
rect 2044 11936 2060 12000
rect 2124 11936 2140 12000
rect 2204 11936 2220 12000
rect 2284 11996 7740 12000
rect 2332 11940 2356 11996
rect 2412 11940 5485 11996
rect 5541 11940 7740 11996
rect 2284 11936 7740 11940
rect 7804 11936 7820 12000
rect 7884 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8220 12000
rect 8284 11996 13740 12000
rect 8284 11940 8375 11996
rect 8431 11940 11265 11996
rect 11321 11940 13740 11996
rect 8284 11936 13740 11940
rect 13804 11936 13820 12000
rect 13884 11936 13900 12000
rect 13964 11936 13980 12000
rect 14044 11936 14060 12000
rect 14124 11936 14140 12000
rect 14204 11996 14220 12000
rect 14211 11940 14220 11996
rect 14204 11936 14220 11940
rect 14284 11996 19740 12000
rect 14284 11940 17045 11996
rect 17101 11940 19740 11996
rect 14284 11936 19740 11940
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11996 19980 12000
rect 19964 11936 19980 11940
rect 20044 11936 20060 12000
rect 20124 11936 20140 12000
rect 20204 11936 20220 12000
rect 20284 11996 25740 12000
rect 20284 11940 22825 11996
rect 22881 11940 25715 11996
rect 20284 11936 25740 11940
rect 25804 11936 25820 12000
rect 25884 11936 25900 12000
rect 25964 11936 25980 12000
rect 26044 11936 26060 12000
rect 26124 11936 26140 12000
rect 26204 11936 26220 12000
rect 26284 11996 31740 12000
rect 26284 11940 28605 11996
rect 28661 11940 31495 11996
rect 31551 11940 31740 11996
rect 26284 11936 31740 11940
rect 31804 11936 31820 12000
rect 31884 11936 31900 12000
rect 31964 11936 31980 12000
rect 32044 11936 32060 12000
rect 32124 11936 32140 12000
rect 32204 11936 32220 12000
rect 32284 11996 37740 12000
rect 32284 11940 34385 11996
rect 34441 11940 37275 11996
rect 37331 11940 37740 11996
rect 32284 11936 37740 11940
rect 37804 11936 37820 12000
rect 37884 11936 37900 12000
rect 37964 11936 37980 12000
rect 38044 11936 38060 12000
rect 38124 11936 38140 12000
rect 38204 11936 38220 12000
rect 38284 11996 43740 12000
rect 38284 11940 40165 11996
rect 40221 11940 43055 11996
rect 43111 11940 43740 11996
rect 38284 11936 43740 11940
rect 43804 11936 43820 12000
rect 43884 11936 43900 12000
rect 43964 11936 43980 12000
rect 44044 11936 44060 12000
rect 44124 11936 44140 12000
rect 44204 11936 44220 12000
rect 44284 11996 49740 12000
rect 49804 11996 49820 12000
rect 49884 11996 49900 12000
rect 44284 11940 45945 11996
rect 46001 11940 48892 11996
rect 48948 11940 49740 11996
rect 49810 11940 49820 11996
rect 49890 11940 49900 11996
rect 44284 11936 49740 11940
rect 49804 11936 49820 11940
rect 49884 11936 49900 11940
rect 49964 11936 49980 12000
rect 50044 11936 50060 12000
rect 50124 11936 50140 12000
rect 50204 11936 50220 12000
rect 50284 11996 55740 12000
rect 50284 11940 53048 11996
rect 53104 11940 53206 11996
rect 53262 11940 53562 11996
rect 53618 11940 54880 11996
rect 54936 11940 55473 11996
rect 55529 11940 55740 11996
rect 50284 11936 55740 11940
rect 55804 11936 55820 12000
rect 55884 11936 55900 12000
rect 55964 11936 55980 12000
rect 56044 11936 56060 12000
rect 56124 11936 56140 12000
rect 56204 11936 56220 12000
rect 56284 11996 61740 12000
rect 56284 11940 56619 11996
rect 56675 11940 58055 11996
rect 58111 11940 58135 11996
rect 58191 11940 59298 11996
rect 59354 11940 59456 11996
rect 59512 11940 59764 11996
rect 59820 11940 59910 11996
rect 59966 11940 60046 11996
rect 60102 11940 60126 11996
rect 60182 11940 61740 11996
rect 56284 11936 61740 11940
rect 61804 11936 61820 12000
rect 61884 11936 61900 12000
rect 61964 11936 61980 12000
rect 62044 11936 62060 12000
rect 62124 11936 62140 12000
rect 62204 11936 62220 12000
rect 62284 11996 67740 12000
rect 62284 11940 62418 11996
rect 62474 11940 62498 11996
rect 62554 11940 67740 11996
rect 62284 11936 67740 11940
rect 67804 11936 67820 12000
rect 67884 11936 67900 12000
rect 67964 11936 67980 12000
rect 68044 11936 68060 12000
rect 68124 11936 68140 12000
rect 68204 11936 68220 12000
rect 68284 11996 73740 12000
rect 68284 11940 71864 11996
rect 71920 11940 71944 11996
rect 72000 11940 72024 11996
rect 72080 11940 72104 11996
rect 72160 11940 73740 11996
rect 68284 11936 73740 11940
rect 73804 11936 73820 12000
rect 73884 11936 73900 12000
rect 73964 11936 73980 12000
rect 74044 11936 74060 12000
rect 74124 11936 74140 12000
rect 74204 11936 74220 12000
rect 74284 11936 75028 12000
rect 964 11912 75028 11936
rect 64454 11732 64460 11796
rect 64524 11794 64530 11796
rect 64597 11794 64663 11797
rect 64524 11792 64663 11794
rect 64524 11736 64602 11792
rect 64658 11736 64663 11792
rect 64524 11734 64663 11736
rect 64524 11732 64530 11734
rect 64597 11731 64663 11734
rect 65333 11794 65399 11797
rect 65926 11794 65932 11796
rect 65333 11792 65932 11794
rect 65333 11736 65338 11792
rect 65394 11736 65932 11792
rect 65333 11734 65932 11736
rect 65333 11731 65399 11734
rect 65926 11732 65932 11734
rect 65996 11732 66002 11796
rect 63350 11460 63356 11524
rect 63420 11522 63426 11524
rect 63585 11522 63651 11525
rect 63420 11520 63651 11522
rect 63420 11464 63590 11520
rect 63646 11464 63651 11520
rect 63420 11462 63651 11464
rect 63420 11460 63426 11462
rect 63585 11459 63651 11462
rect 62982 10508 62988 10572
rect 63052 10570 63058 10572
rect 63585 10570 63651 10573
rect 63052 10568 63651 10570
rect 63052 10512 63590 10568
rect 63646 10512 63651 10568
rect 63052 10510 63651 10512
rect 63052 10508 63058 10510
rect 63585 10507 63651 10510
rect 63350 9964 63356 10028
rect 63420 10026 63426 10028
rect 63493 10026 63559 10029
rect 63420 10024 63559 10026
rect 63420 9968 63498 10024
rect 63554 9968 63559 10024
rect 63420 9966 63559 9968
rect 63420 9964 63426 9966
rect 63493 9963 63559 9966
rect 63166 9828 63172 9892
rect 63236 9890 63242 9892
rect 63493 9890 63559 9893
rect 63236 9888 63559 9890
rect 63236 9832 63498 9888
rect 63554 9832 63559 9888
rect 63236 9830 63559 9832
rect 63236 9828 63242 9830
rect 63493 9827 63559 9830
rect 66069 9210 66135 9213
rect 66069 9208 66178 9210
rect 66069 9152 66074 9208
rect 66130 9152 66178 9208
rect 66069 9147 66178 9152
rect 66118 8941 66178 9147
rect 66118 8936 66227 8941
rect 66118 8880 66166 8936
rect 66222 8880 66227 8936
rect 66118 8878 66227 8880
rect 66161 8875 66227 8878
rect 59269 7850 59335 7853
rect 65742 7850 65748 7852
rect 59269 7848 65748 7850
rect 59269 7792 59274 7848
rect 59330 7792 65748 7848
rect 59269 7790 65748 7792
rect 59269 7787 59335 7790
rect 65742 7788 65748 7790
rect 65812 7788 65818 7852
rect 66253 7850 66319 7853
rect 66253 7848 66362 7850
rect 66253 7792 66258 7848
rect 66314 7792 66362 7848
rect 66253 7787 66362 7792
rect 59629 7714 59695 7717
rect 61285 7714 61351 7717
rect 59629 7712 61351 7714
rect 59629 7656 59634 7712
rect 59690 7656 61290 7712
rect 61346 7656 61351 7712
rect 59629 7654 61351 7656
rect 59629 7651 59695 7654
rect 61285 7651 61351 7654
rect 61469 7714 61535 7717
rect 64597 7714 64663 7717
rect 61469 7712 64663 7714
rect 61469 7656 61474 7712
rect 61530 7656 64602 7712
rect 64658 7656 64663 7712
rect 61469 7654 64663 7656
rect 61469 7651 61535 7654
rect 64597 7651 64663 7654
rect 58249 7578 58315 7581
rect 63534 7578 63540 7580
rect 58249 7576 63540 7578
rect 58249 7520 58254 7576
rect 58310 7520 63540 7576
rect 58249 7518 63540 7520
rect 58249 7515 58315 7518
rect 63534 7516 63540 7518
rect 63604 7516 63610 7580
rect 61285 7442 61351 7445
rect 66110 7442 66116 7444
rect 61285 7440 66116 7442
rect 61285 7384 61290 7440
rect 61346 7384 66116 7440
rect 61285 7382 66116 7384
rect 61285 7379 61351 7382
rect 66110 7380 66116 7382
rect 66180 7380 66186 7444
rect 66302 7442 66362 7787
rect 66437 7442 66503 7445
rect 66302 7440 66503 7442
rect 66302 7384 66442 7440
rect 66498 7384 66503 7440
rect 66302 7382 66503 7384
rect 66437 7379 66503 7382
rect 62665 7306 62731 7309
rect 67030 7306 67036 7308
rect 62665 7304 67036 7306
rect 62665 7248 62670 7304
rect 62726 7248 67036 7304
rect 62665 7246 67036 7248
rect 62665 7243 62731 7246
rect 67030 7244 67036 7246
rect 67100 7244 67106 7308
rect 57329 7170 57395 7173
rect 62982 7170 62988 7172
rect 57329 7168 62988 7170
rect 57329 7112 57334 7168
rect 57390 7112 62988 7168
rect 57329 7110 62988 7112
rect 57329 7107 57395 7110
rect 62982 7108 62988 7110
rect 63052 7108 63058 7172
rect 62573 7034 62639 7037
rect 66294 7034 66300 7036
rect 62573 7032 66300 7034
rect 62573 6976 62578 7032
rect 62634 6976 66300 7032
rect 62573 6974 66300 6976
rect 62573 6971 62639 6974
rect 66294 6972 66300 6974
rect 66364 6972 66370 7036
rect 55029 6762 55095 6765
rect 63902 6762 63908 6764
rect 55029 6760 63908 6762
rect 55029 6704 55034 6760
rect 55090 6704 63908 6760
rect 55029 6702 63908 6704
rect 55029 6699 55095 6702
rect 63902 6700 63908 6702
rect 63972 6700 63978 6764
rect 52361 6626 52427 6629
rect 64270 6626 64276 6628
rect 52361 6624 64276 6626
rect 52361 6568 52366 6624
rect 52422 6568 64276 6624
rect 52361 6566 64276 6568
rect 52361 6563 52427 6566
rect 64270 6564 64276 6566
rect 64340 6564 64346 6628
rect 40217 6490 40283 6493
rect 64321 6490 64387 6493
rect 40217 6488 64387 6490
rect 40217 6432 40222 6488
rect 40278 6432 64326 6488
rect 64382 6432 64387 6488
rect 40217 6430 64387 6432
rect 40217 6427 40283 6430
rect 64321 6427 64387 6430
rect 33777 6354 33843 6357
rect 67817 6354 67883 6357
rect 33777 6352 67883 6354
rect 33777 6296 33782 6352
rect 33838 6296 67822 6352
rect 67878 6296 67883 6352
rect 33777 6294 67883 6296
rect 33777 6291 33843 6294
rect 67817 6291 67883 6294
rect 31569 6218 31635 6221
rect 67633 6218 67699 6221
rect 31569 6216 67699 6218
rect 31569 6160 31574 6216
rect 31630 6160 67638 6216
rect 67694 6160 67699 6216
rect 31569 6158 67699 6160
rect 31569 6155 31635 6158
rect 67633 6155 67699 6158
rect 62849 6082 62915 6085
rect 63585 6082 63651 6085
rect 62849 6080 63651 6082
rect 62849 6024 62854 6080
rect 62910 6024 63590 6080
rect 63646 6024 63651 6080
rect 62849 6022 63651 6024
rect 62849 6019 62915 6022
rect 63585 6019 63651 6022
rect 56501 5946 56567 5949
rect 63718 5946 63724 5948
rect 56501 5944 63724 5946
rect 56501 5888 56506 5944
rect 56562 5888 63724 5944
rect 56501 5886 63724 5888
rect 56501 5883 56567 5886
rect 63718 5884 63724 5886
rect 63788 5884 63794 5948
rect 44725 5810 44791 5813
rect 69473 5810 69539 5813
rect 44725 5808 69539 5810
rect 44725 5752 44730 5808
rect 44786 5752 69478 5808
rect 69534 5752 69539 5808
rect 44725 5750 69539 5752
rect 44725 5747 44791 5750
rect 69473 5747 69539 5750
rect 42701 5674 42767 5677
rect 68553 5674 68619 5677
rect 42701 5672 68619 5674
rect 42701 5616 42706 5672
rect 42762 5616 68558 5672
rect 68614 5616 68619 5672
rect 42701 5614 68619 5616
rect 42701 5611 42767 5614
rect 68553 5611 68619 5614
rect 53741 5538 53807 5541
rect 63350 5538 63356 5540
rect 53741 5536 63356 5538
rect 53741 5480 53746 5536
rect 53802 5480 63356 5536
rect 53741 5478 63356 5480
rect 53741 5475 53807 5478
rect 63350 5476 63356 5478
rect 63420 5476 63426 5540
rect 30741 5402 30807 5405
rect 34881 5402 34947 5405
rect 35801 5402 35867 5405
rect 30741 5400 35867 5402
rect 30741 5344 30746 5400
rect 30802 5344 34886 5400
rect 34942 5344 35806 5400
rect 35862 5344 35867 5400
rect 30741 5342 35867 5344
rect 30741 5339 30807 5342
rect 34881 5339 34947 5342
rect 35801 5339 35867 5342
rect 31661 5266 31727 5269
rect 32213 5266 32279 5269
rect 31661 5264 32279 5266
rect 31661 5208 31666 5264
rect 31722 5208 32218 5264
rect 32274 5208 32279 5264
rect 31661 5206 32279 5208
rect 31661 5203 31727 5206
rect 32213 5203 32279 5206
rect 32489 5266 32555 5269
rect 37917 5266 37983 5269
rect 32489 5264 37983 5266
rect 32489 5208 32494 5264
rect 32550 5208 37922 5264
rect 37978 5208 37983 5264
rect 32489 5206 37983 5208
rect 32489 5203 32555 5206
rect 37917 5203 37983 5206
rect 61745 5266 61811 5269
rect 62389 5266 62455 5269
rect 61745 5264 62455 5266
rect 61745 5208 61750 5264
rect 61806 5208 62394 5264
rect 62450 5208 62455 5264
rect 61745 5206 62455 5208
rect 61745 5203 61811 5206
rect 62389 5203 62455 5206
rect 30925 5130 30991 5133
rect 32397 5130 32463 5133
rect 30925 5128 32463 5130
rect 30925 5072 30930 5128
rect 30986 5072 32402 5128
rect 32458 5072 32463 5128
rect 30925 5070 32463 5072
rect 30925 5067 30991 5070
rect 32397 5067 32463 5070
rect 34053 5130 34119 5133
rect 35617 5130 35683 5133
rect 34053 5128 35683 5130
rect 34053 5072 34058 5128
rect 34114 5072 35622 5128
rect 35678 5072 35683 5128
rect 34053 5070 35683 5072
rect 34053 5067 34119 5070
rect 35617 5067 35683 5070
rect 60273 5130 60339 5133
rect 65241 5130 65307 5133
rect 60273 5128 65307 5130
rect 60273 5072 60278 5128
rect 60334 5072 65246 5128
rect 65302 5072 65307 5128
rect 60273 5070 65307 5072
rect 60273 5067 60339 5070
rect 65241 5067 65307 5070
rect 32397 4994 32463 4997
rect 36261 4994 36327 4997
rect 32397 4992 36327 4994
rect 32397 4936 32402 4992
rect 32458 4936 36266 4992
rect 36322 4936 36327 4992
rect 32397 4934 36327 4936
rect 32397 4931 32463 4934
rect 36261 4931 36327 4934
rect 45277 4994 45343 4997
rect 48497 4994 48563 4997
rect 45277 4992 48563 4994
rect 45277 4936 45282 4992
rect 45338 4936 48502 4992
rect 48558 4936 48563 4992
rect 45277 4934 48563 4936
rect 45277 4931 45343 4934
rect 48497 4931 48563 4934
rect 60457 4994 60523 4997
rect 61101 4994 61167 4997
rect 60457 4992 61167 4994
rect 60457 4936 60462 4992
rect 60518 4936 61106 4992
rect 61162 4936 61167 4992
rect 60457 4934 61167 4936
rect 60457 4931 60523 4934
rect 61101 4931 61167 4934
rect 33961 4860 34027 4861
rect 33910 4858 33916 4860
rect 33870 4798 33916 4858
rect 33980 4856 34027 4860
rect 34022 4800 34027 4856
rect 33910 4796 33916 4798
rect 33980 4796 34027 4800
rect 33961 4795 34027 4796
rect 34697 4858 34763 4861
rect 34973 4858 35039 4861
rect 68645 4858 68711 4861
rect 34697 4856 68711 4858
rect 34697 4800 34702 4856
rect 34758 4800 34978 4856
rect 35034 4800 68650 4856
rect 68706 4800 68711 4856
rect 34697 4798 68711 4800
rect 34697 4795 34763 4798
rect 34973 4795 35039 4798
rect 68645 4795 68711 4798
rect 964 4592 75028 4616
rect 964 4588 4740 4592
rect 964 4532 4216 4588
rect 4272 4532 4296 4588
rect 4352 4532 4376 4588
rect 4432 4532 4456 4588
rect 4512 4532 4740 4588
rect 964 4528 4740 4532
rect 4804 4528 4820 4592
rect 4884 4528 4900 4592
rect 4964 4528 4980 4592
rect 5044 4528 5060 4592
rect 5124 4528 5140 4592
rect 5204 4528 5220 4592
rect 5284 4528 10740 4592
rect 10804 4528 10820 4592
rect 10884 4528 10900 4592
rect 10964 4528 10980 4592
rect 11044 4528 11060 4592
rect 11124 4528 11140 4592
rect 11204 4528 11220 4592
rect 11284 4588 16740 4592
rect 11284 4532 14216 4588
rect 14272 4532 14296 4588
rect 14352 4532 14376 4588
rect 14432 4532 14456 4588
rect 14512 4532 16740 4588
rect 11284 4528 16740 4532
rect 16804 4528 16820 4592
rect 16884 4528 16900 4592
rect 16964 4528 16980 4592
rect 17044 4528 17060 4592
rect 17124 4528 17140 4592
rect 17204 4528 17220 4592
rect 17284 4528 22740 4592
rect 22804 4528 22820 4592
rect 22884 4528 22900 4592
rect 22964 4528 22980 4592
rect 23044 4528 23060 4592
rect 23124 4528 23140 4592
rect 23204 4528 23220 4592
rect 23284 4588 28740 4592
rect 23284 4532 24216 4588
rect 24272 4532 24296 4588
rect 24352 4532 24376 4588
rect 24432 4532 24456 4588
rect 24512 4532 28740 4588
rect 23284 4528 28740 4532
rect 28804 4528 28820 4592
rect 28884 4528 28900 4592
rect 28964 4528 28980 4592
rect 29044 4528 29060 4592
rect 29124 4528 29140 4592
rect 29204 4528 29220 4592
rect 29284 4588 34740 4592
rect 29284 4532 34216 4588
rect 34272 4532 34296 4588
rect 34352 4532 34376 4588
rect 34432 4532 34456 4588
rect 34512 4532 34740 4588
rect 29284 4528 34740 4532
rect 34804 4528 34820 4592
rect 34884 4528 34900 4592
rect 34964 4528 34980 4592
rect 35044 4528 35060 4592
rect 35124 4528 35140 4592
rect 35204 4528 35220 4592
rect 35284 4528 40740 4592
rect 40804 4528 40820 4592
rect 40884 4528 40900 4592
rect 40964 4528 40980 4592
rect 41044 4528 41060 4592
rect 41124 4528 41140 4592
rect 41204 4528 41220 4592
rect 41284 4588 46740 4592
rect 41284 4532 44216 4588
rect 44272 4532 44296 4588
rect 44352 4532 44376 4588
rect 44432 4532 44456 4588
rect 44512 4532 46740 4588
rect 41284 4528 46740 4532
rect 46804 4528 46820 4592
rect 46884 4528 46900 4592
rect 46964 4528 46980 4592
rect 47044 4528 47060 4592
rect 47124 4528 47140 4592
rect 47204 4528 47220 4592
rect 47284 4528 52740 4592
rect 52804 4528 52820 4592
rect 52884 4528 52900 4592
rect 52964 4528 52980 4592
rect 53044 4528 53060 4592
rect 53124 4528 53140 4592
rect 53204 4528 53220 4592
rect 53284 4588 58740 4592
rect 53284 4532 54216 4588
rect 54272 4532 54296 4588
rect 54352 4532 54376 4588
rect 54432 4532 54456 4588
rect 54512 4532 58740 4588
rect 53284 4528 58740 4532
rect 58804 4528 58820 4592
rect 58884 4528 58900 4592
rect 58964 4528 58980 4592
rect 59044 4528 59060 4592
rect 59124 4528 59140 4592
rect 59204 4528 59220 4592
rect 59284 4588 64740 4592
rect 59284 4532 64216 4588
rect 64272 4532 64296 4588
rect 64352 4532 64376 4588
rect 64432 4532 64456 4588
rect 64512 4532 64740 4588
rect 59284 4528 64740 4532
rect 64804 4528 64820 4592
rect 64884 4528 64900 4592
rect 64964 4528 64980 4592
rect 65044 4528 65060 4592
rect 65124 4528 65140 4592
rect 65204 4528 65220 4592
rect 65284 4528 70740 4592
rect 70804 4528 70820 4592
rect 70884 4528 70900 4592
rect 70964 4528 70980 4592
rect 71044 4528 71060 4592
rect 71124 4528 71140 4592
rect 71204 4528 71220 4592
rect 71284 4588 75028 4592
rect 71284 4532 74216 4588
rect 74272 4532 74296 4588
rect 74352 4532 74376 4588
rect 74432 4532 74456 4588
rect 74512 4532 75028 4588
rect 71284 4528 75028 4532
rect 964 4512 75028 4528
rect 964 4508 4740 4512
rect 964 4452 4216 4508
rect 4272 4452 4296 4508
rect 4352 4452 4376 4508
rect 4432 4452 4456 4508
rect 4512 4452 4740 4508
rect 964 4448 4740 4452
rect 4804 4448 4820 4512
rect 4884 4448 4900 4512
rect 4964 4448 4980 4512
rect 5044 4448 5060 4512
rect 5124 4448 5140 4512
rect 5204 4448 5220 4512
rect 5284 4448 10740 4512
rect 10804 4448 10820 4512
rect 10884 4448 10900 4512
rect 10964 4448 10980 4512
rect 11044 4448 11060 4512
rect 11124 4448 11140 4512
rect 11204 4448 11220 4512
rect 11284 4508 16740 4512
rect 11284 4452 14216 4508
rect 14272 4452 14296 4508
rect 14352 4452 14376 4508
rect 14432 4452 14456 4508
rect 14512 4452 16740 4508
rect 11284 4448 16740 4452
rect 16804 4448 16820 4512
rect 16884 4448 16900 4512
rect 16964 4448 16980 4512
rect 17044 4448 17060 4512
rect 17124 4448 17140 4512
rect 17204 4448 17220 4512
rect 17284 4448 22740 4512
rect 22804 4448 22820 4512
rect 22884 4448 22900 4512
rect 22964 4448 22980 4512
rect 23044 4448 23060 4512
rect 23124 4448 23140 4512
rect 23204 4448 23220 4512
rect 23284 4508 28740 4512
rect 23284 4452 24216 4508
rect 24272 4452 24296 4508
rect 24352 4452 24376 4508
rect 24432 4452 24456 4508
rect 24512 4452 28740 4508
rect 23284 4448 28740 4452
rect 28804 4448 28820 4512
rect 28884 4448 28900 4512
rect 28964 4448 28980 4512
rect 29044 4448 29060 4512
rect 29124 4448 29140 4512
rect 29204 4448 29220 4512
rect 29284 4508 34740 4512
rect 29284 4452 34216 4508
rect 34272 4452 34296 4508
rect 34352 4452 34376 4508
rect 34432 4452 34456 4508
rect 34512 4452 34740 4508
rect 29284 4448 34740 4452
rect 34804 4448 34820 4512
rect 34884 4448 34900 4512
rect 34964 4448 34980 4512
rect 35044 4448 35060 4512
rect 35124 4448 35140 4512
rect 35204 4448 35220 4512
rect 35284 4448 40740 4512
rect 40804 4448 40820 4512
rect 40884 4448 40900 4512
rect 40964 4448 40980 4512
rect 41044 4448 41060 4512
rect 41124 4448 41140 4512
rect 41204 4448 41220 4512
rect 41284 4508 46740 4512
rect 41284 4452 44216 4508
rect 44272 4452 44296 4508
rect 44352 4452 44376 4508
rect 44432 4452 44456 4508
rect 44512 4452 46740 4508
rect 41284 4448 46740 4452
rect 46804 4448 46820 4512
rect 46884 4448 46900 4512
rect 46964 4448 46980 4512
rect 47044 4448 47060 4512
rect 47124 4448 47140 4512
rect 47204 4448 47220 4512
rect 47284 4448 52740 4512
rect 52804 4448 52820 4512
rect 52884 4448 52900 4512
rect 52964 4448 52980 4512
rect 53044 4448 53060 4512
rect 53124 4448 53140 4512
rect 53204 4448 53220 4512
rect 53284 4508 58740 4512
rect 53284 4452 54216 4508
rect 54272 4452 54296 4508
rect 54352 4452 54376 4508
rect 54432 4452 54456 4508
rect 54512 4452 58740 4508
rect 53284 4448 58740 4452
rect 58804 4448 58820 4512
rect 58884 4448 58900 4512
rect 58964 4448 58980 4512
rect 59044 4448 59060 4512
rect 59124 4448 59140 4512
rect 59204 4448 59220 4512
rect 59284 4508 64740 4512
rect 59284 4452 64216 4508
rect 64272 4452 64296 4508
rect 64352 4452 64376 4508
rect 64432 4452 64456 4508
rect 64512 4452 64740 4508
rect 59284 4448 64740 4452
rect 64804 4448 64820 4512
rect 64884 4448 64900 4512
rect 64964 4448 64980 4512
rect 65044 4448 65060 4512
rect 65124 4448 65140 4512
rect 65204 4448 65220 4512
rect 65284 4448 70740 4512
rect 70804 4448 70820 4512
rect 70884 4448 70900 4512
rect 70964 4448 70980 4512
rect 71044 4448 71060 4512
rect 71124 4448 71140 4512
rect 71204 4448 71220 4512
rect 71284 4508 75028 4512
rect 71284 4452 74216 4508
rect 74272 4452 74296 4508
rect 74352 4452 74376 4508
rect 74432 4452 74456 4508
rect 74512 4452 75028 4508
rect 71284 4448 75028 4452
rect 964 4432 75028 4448
rect 964 4428 4740 4432
rect 964 4372 4216 4428
rect 4272 4372 4296 4428
rect 4352 4372 4376 4428
rect 4432 4372 4456 4428
rect 4512 4372 4740 4428
rect 964 4368 4740 4372
rect 4804 4368 4820 4432
rect 4884 4368 4900 4432
rect 4964 4368 4980 4432
rect 5044 4368 5060 4432
rect 5124 4368 5140 4432
rect 5204 4368 5220 4432
rect 5284 4368 10740 4432
rect 10804 4368 10820 4432
rect 10884 4368 10900 4432
rect 10964 4368 10980 4432
rect 11044 4368 11060 4432
rect 11124 4368 11140 4432
rect 11204 4368 11220 4432
rect 11284 4428 16740 4432
rect 11284 4372 14216 4428
rect 14272 4372 14296 4428
rect 14352 4372 14376 4428
rect 14432 4372 14456 4428
rect 14512 4372 16740 4428
rect 11284 4368 16740 4372
rect 16804 4368 16820 4432
rect 16884 4368 16900 4432
rect 16964 4368 16980 4432
rect 17044 4368 17060 4432
rect 17124 4368 17140 4432
rect 17204 4368 17220 4432
rect 17284 4368 22740 4432
rect 22804 4368 22820 4432
rect 22884 4368 22900 4432
rect 22964 4368 22980 4432
rect 23044 4368 23060 4432
rect 23124 4368 23140 4432
rect 23204 4368 23220 4432
rect 23284 4428 28740 4432
rect 23284 4372 24216 4428
rect 24272 4372 24296 4428
rect 24352 4372 24376 4428
rect 24432 4372 24456 4428
rect 24512 4372 28740 4428
rect 23284 4368 28740 4372
rect 28804 4368 28820 4432
rect 28884 4368 28900 4432
rect 28964 4368 28980 4432
rect 29044 4368 29060 4432
rect 29124 4368 29140 4432
rect 29204 4368 29220 4432
rect 29284 4428 34740 4432
rect 29284 4372 34216 4428
rect 34272 4372 34296 4428
rect 34352 4372 34376 4428
rect 34432 4372 34456 4428
rect 34512 4372 34740 4428
rect 29284 4368 34740 4372
rect 34804 4368 34820 4432
rect 34884 4368 34900 4432
rect 34964 4368 34980 4432
rect 35044 4368 35060 4432
rect 35124 4368 35140 4432
rect 35204 4368 35220 4432
rect 35284 4368 40740 4432
rect 40804 4368 40820 4432
rect 40884 4368 40900 4432
rect 40964 4368 40980 4432
rect 41044 4368 41060 4432
rect 41124 4368 41140 4432
rect 41204 4368 41220 4432
rect 41284 4428 46740 4432
rect 41284 4372 44216 4428
rect 44272 4372 44296 4428
rect 44352 4372 44376 4428
rect 44432 4372 44456 4428
rect 44512 4372 46740 4428
rect 41284 4368 46740 4372
rect 46804 4368 46820 4432
rect 46884 4368 46900 4432
rect 46964 4368 46980 4432
rect 47044 4368 47060 4432
rect 47124 4368 47140 4432
rect 47204 4368 47220 4432
rect 47284 4368 52740 4432
rect 52804 4368 52820 4432
rect 52884 4368 52900 4432
rect 52964 4368 52980 4432
rect 53044 4368 53060 4432
rect 53124 4368 53140 4432
rect 53204 4368 53220 4432
rect 53284 4428 58740 4432
rect 53284 4372 54216 4428
rect 54272 4372 54296 4428
rect 54352 4372 54376 4428
rect 54432 4372 54456 4428
rect 54512 4372 58740 4428
rect 53284 4368 58740 4372
rect 58804 4368 58820 4432
rect 58884 4368 58900 4432
rect 58964 4368 58980 4432
rect 59044 4368 59060 4432
rect 59124 4368 59140 4432
rect 59204 4368 59220 4432
rect 59284 4428 64740 4432
rect 59284 4372 64216 4428
rect 64272 4372 64296 4428
rect 64352 4372 64376 4428
rect 64432 4372 64456 4428
rect 64512 4372 64740 4428
rect 59284 4368 64740 4372
rect 64804 4368 64820 4432
rect 64884 4368 64900 4432
rect 64964 4368 64980 4432
rect 65044 4368 65060 4432
rect 65124 4368 65140 4432
rect 65204 4368 65220 4432
rect 65284 4368 70740 4432
rect 70804 4368 70820 4432
rect 70884 4368 70900 4432
rect 70964 4368 70980 4432
rect 71044 4368 71060 4432
rect 71124 4368 71140 4432
rect 71204 4368 71220 4432
rect 71284 4428 75028 4432
rect 71284 4372 74216 4428
rect 74272 4372 74296 4428
rect 74352 4372 74376 4428
rect 74432 4372 74456 4428
rect 74512 4372 75028 4428
rect 71284 4368 75028 4372
rect 964 4352 75028 4368
rect 964 4348 4740 4352
rect 964 4292 4216 4348
rect 4272 4292 4296 4348
rect 4352 4292 4376 4348
rect 4432 4292 4456 4348
rect 4512 4292 4740 4348
rect 964 4288 4740 4292
rect 4804 4288 4820 4352
rect 4884 4288 4900 4352
rect 4964 4288 4980 4352
rect 5044 4288 5060 4352
rect 5124 4288 5140 4352
rect 5204 4288 5220 4352
rect 5284 4288 10740 4352
rect 10804 4288 10820 4352
rect 10884 4288 10900 4352
rect 10964 4288 10980 4352
rect 11044 4288 11060 4352
rect 11124 4288 11140 4352
rect 11204 4288 11220 4352
rect 11284 4348 16740 4352
rect 11284 4292 14216 4348
rect 14272 4292 14296 4348
rect 14352 4292 14376 4348
rect 14432 4292 14456 4348
rect 14512 4292 16740 4348
rect 11284 4288 16740 4292
rect 16804 4288 16820 4352
rect 16884 4288 16900 4352
rect 16964 4288 16980 4352
rect 17044 4288 17060 4352
rect 17124 4288 17140 4352
rect 17204 4288 17220 4352
rect 17284 4288 22740 4352
rect 22804 4288 22820 4352
rect 22884 4288 22900 4352
rect 22964 4288 22980 4352
rect 23044 4288 23060 4352
rect 23124 4288 23140 4352
rect 23204 4288 23220 4352
rect 23284 4348 28740 4352
rect 23284 4292 24216 4348
rect 24272 4292 24296 4348
rect 24352 4292 24376 4348
rect 24432 4292 24456 4348
rect 24512 4292 28740 4348
rect 23284 4288 28740 4292
rect 28804 4288 28820 4352
rect 28884 4288 28900 4352
rect 28964 4288 28980 4352
rect 29044 4288 29060 4352
rect 29124 4288 29140 4352
rect 29204 4288 29220 4352
rect 29284 4348 34740 4352
rect 29284 4292 34216 4348
rect 34272 4292 34296 4348
rect 34352 4292 34376 4348
rect 34432 4292 34456 4348
rect 34512 4292 34740 4348
rect 29284 4288 34740 4292
rect 34804 4288 34820 4352
rect 34884 4288 34900 4352
rect 34964 4288 34980 4352
rect 35044 4288 35060 4352
rect 35124 4288 35140 4352
rect 35204 4288 35220 4352
rect 35284 4288 40740 4352
rect 40804 4288 40820 4352
rect 40884 4288 40900 4352
rect 40964 4288 40980 4352
rect 41044 4288 41060 4352
rect 41124 4288 41140 4352
rect 41204 4288 41220 4352
rect 41284 4348 46740 4352
rect 41284 4292 44216 4348
rect 44272 4292 44296 4348
rect 44352 4292 44376 4348
rect 44432 4292 44456 4348
rect 44512 4292 46740 4348
rect 41284 4288 46740 4292
rect 46804 4288 46820 4352
rect 46884 4288 46900 4352
rect 46964 4288 46980 4352
rect 47044 4288 47060 4352
rect 47124 4288 47140 4352
rect 47204 4288 47220 4352
rect 47284 4288 52740 4352
rect 52804 4288 52820 4352
rect 52884 4288 52900 4352
rect 52964 4288 52980 4352
rect 53044 4288 53060 4352
rect 53124 4288 53140 4352
rect 53204 4288 53220 4352
rect 53284 4348 58740 4352
rect 53284 4292 54216 4348
rect 54272 4292 54296 4348
rect 54352 4292 54376 4348
rect 54432 4292 54456 4348
rect 54512 4292 58740 4348
rect 53284 4288 58740 4292
rect 58804 4288 58820 4352
rect 58884 4288 58900 4352
rect 58964 4288 58980 4352
rect 59044 4288 59060 4352
rect 59124 4288 59140 4352
rect 59204 4288 59220 4352
rect 59284 4348 64740 4352
rect 59284 4292 64216 4348
rect 64272 4292 64296 4348
rect 64352 4292 64376 4348
rect 64432 4292 64456 4348
rect 64512 4292 64740 4348
rect 59284 4288 64740 4292
rect 64804 4288 64820 4352
rect 64884 4288 64900 4352
rect 64964 4288 64980 4352
rect 65044 4288 65060 4352
rect 65124 4288 65140 4352
rect 65204 4288 65220 4352
rect 65284 4288 70740 4352
rect 70804 4288 70820 4352
rect 70884 4288 70900 4352
rect 70964 4288 70980 4352
rect 71044 4288 71060 4352
rect 71124 4288 71140 4352
rect 71204 4288 71220 4352
rect 71284 4348 75028 4352
rect 71284 4292 74216 4348
rect 74272 4292 74296 4348
rect 74352 4292 74376 4348
rect 74432 4292 74456 4348
rect 74512 4292 75028 4348
rect 71284 4288 75028 4292
rect 964 4264 75028 4288
rect 32305 4178 32371 4181
rect 33593 4178 33659 4181
rect 34053 4178 34119 4181
rect 35157 4178 35223 4181
rect 35433 4178 35499 4181
rect 32305 4176 35499 4178
rect 32305 4120 32310 4176
rect 32366 4120 33598 4176
rect 33654 4120 34058 4176
rect 34114 4120 35162 4176
rect 35218 4120 35438 4176
rect 35494 4120 35499 4176
rect 32305 4118 35499 4120
rect 32305 4115 32371 4118
rect 33593 4115 33659 4118
rect 34053 4115 34119 4118
rect 35157 4115 35223 4118
rect 35433 4115 35499 4118
rect 61193 4178 61259 4181
rect 63677 4178 63743 4181
rect 61193 4176 63743 4178
rect 61193 4120 61198 4176
rect 61254 4120 63682 4176
rect 63738 4120 63743 4176
rect 61193 4118 63743 4120
rect 61193 4115 61259 4118
rect 63677 4115 63743 4118
rect 29821 4042 29887 4045
rect 65793 4042 65859 4045
rect 29821 4040 65859 4042
rect 29821 3984 29826 4040
rect 29882 3984 65798 4040
rect 65854 3984 65859 4040
rect 29821 3982 65859 3984
rect 29821 3979 29887 3982
rect 65793 3979 65859 3982
rect 33409 3906 33475 3909
rect 36261 3906 36327 3909
rect 66478 3906 66484 3908
rect 33409 3904 36186 3906
rect 33409 3848 33414 3904
rect 33470 3848 36186 3904
rect 33409 3846 36186 3848
rect 33409 3843 33475 3846
rect 33961 3770 34027 3773
rect 35249 3770 35315 3773
rect 35709 3770 35775 3773
rect 33961 3768 35775 3770
rect 33961 3712 33966 3768
rect 34022 3712 35254 3768
rect 35310 3712 35714 3768
rect 35770 3712 35775 3768
rect 33961 3710 35775 3712
rect 36126 3770 36186 3846
rect 36261 3904 66484 3906
rect 36261 3848 36266 3904
rect 36322 3848 66484 3904
rect 36261 3846 66484 3848
rect 36261 3843 36327 3846
rect 66478 3844 66484 3846
rect 66548 3844 66554 3908
rect 36629 3770 36695 3773
rect 36126 3768 36695 3770
rect 36126 3712 36634 3768
rect 36690 3712 36695 3768
rect 36126 3710 36695 3712
rect 33961 3707 34027 3710
rect 35249 3707 35315 3710
rect 35709 3707 35775 3710
rect 36629 3707 36695 3710
rect 50337 3770 50403 3773
rect 69054 3770 69060 3772
rect 50337 3768 69060 3770
rect 50337 3712 50342 3768
rect 50398 3712 69060 3768
rect 50337 3710 69060 3712
rect 50337 3707 50403 3710
rect 69054 3708 69060 3710
rect 69124 3708 69130 3772
rect 32581 3634 32647 3637
rect 69933 3634 69999 3637
rect 32581 3632 69999 3634
rect 32581 3576 32586 3632
rect 32642 3576 69938 3632
rect 69994 3576 69999 3632
rect 32581 3574 69999 3576
rect 32581 3571 32647 3574
rect 69933 3571 69999 3574
rect 26877 3498 26943 3501
rect 66069 3498 66135 3501
rect 26877 3496 66135 3498
rect 26877 3440 26882 3496
rect 26938 3440 66074 3496
rect 66130 3440 66135 3496
rect 26877 3438 66135 3440
rect 26877 3435 26943 3438
rect 66069 3435 66135 3438
rect 32397 3362 32463 3365
rect 33777 3362 33843 3365
rect 32397 3360 33843 3362
rect 32397 3304 32402 3360
rect 32458 3304 33782 3360
rect 33838 3304 33843 3360
rect 32397 3302 33843 3304
rect 32397 3299 32463 3302
rect 33777 3299 33843 3302
rect 33961 3362 34027 3365
rect 34973 3362 35039 3365
rect 33961 3360 35039 3362
rect 33961 3304 33966 3360
rect 34022 3304 34978 3360
rect 35034 3304 35039 3360
rect 33961 3302 35039 3304
rect 33961 3299 34027 3302
rect 34973 3299 35039 3302
rect 53005 3362 53071 3365
rect 53373 3362 53439 3365
rect 64086 3362 64092 3364
rect 53005 3360 64092 3362
rect 53005 3304 53010 3360
rect 53066 3304 53378 3360
rect 53434 3304 64092 3360
rect 53005 3302 64092 3304
rect 53005 3299 53071 3302
rect 53373 3299 53439 3302
rect 64086 3300 64092 3302
rect 64156 3300 64162 3364
rect 31661 3226 31727 3229
rect 36077 3226 36143 3229
rect 31661 3224 36143 3226
rect 31661 3168 31666 3224
rect 31722 3168 36082 3224
rect 36138 3168 36143 3224
rect 31661 3166 36143 3168
rect 31661 3163 31727 3166
rect 36077 3163 36143 3166
rect 50889 3226 50955 3229
rect 51165 3226 51231 3229
rect 50889 3224 51231 3226
rect 50889 3168 50894 3224
rect 50950 3168 51170 3224
rect 51226 3168 51231 3224
rect 50889 3166 51231 3168
rect 50889 3163 50955 3166
rect 51165 3163 51231 3166
rect 58709 3226 58775 3229
rect 62389 3226 62455 3229
rect 58709 3224 62455 3226
rect 58709 3168 58714 3224
rect 58770 3168 62394 3224
rect 62450 3168 62455 3224
rect 58709 3166 62455 3168
rect 58709 3163 58775 3166
rect 62389 3163 62455 3166
rect 32213 3090 32279 3093
rect 36445 3090 36511 3093
rect 32213 3088 36511 3090
rect 32213 3032 32218 3088
rect 32274 3032 36450 3088
rect 36506 3032 36511 3088
rect 32213 3030 36511 3032
rect 32213 3027 32279 3030
rect 36445 3027 36511 3030
rect 37457 3090 37523 3093
rect 67214 3090 67220 3092
rect 37457 3088 67220 3090
rect 37457 3032 37462 3088
rect 37518 3032 67220 3088
rect 37457 3030 67220 3032
rect 37457 3027 37523 3030
rect 67214 3028 67220 3030
rect 67284 3028 67290 3092
rect 33409 2954 33475 2957
rect 35433 2954 35499 2957
rect 33409 2952 35499 2954
rect 33409 2896 33414 2952
rect 33470 2896 35438 2952
rect 35494 2896 35499 2952
rect 33409 2894 35499 2896
rect 33409 2891 33475 2894
rect 35433 2891 35499 2894
rect 29729 2818 29795 2821
rect 36169 2818 36235 2821
rect 29729 2816 36235 2818
rect 29729 2760 29734 2816
rect 29790 2760 36174 2816
rect 36230 2760 36235 2816
rect 29729 2758 36235 2760
rect 29729 2755 29795 2758
rect 36169 2755 36235 2758
rect 33869 2548 33935 2549
rect 33869 2546 33916 2548
rect 33824 2544 33916 2546
rect 33824 2488 33874 2544
rect 33824 2486 33916 2488
rect 33869 2484 33916 2486
rect 33980 2484 33986 2548
rect 33869 2483 33935 2484
rect 30557 2410 30623 2413
rect 34881 2410 34947 2413
rect 30557 2408 34947 2410
rect 30557 2352 30562 2408
rect 30618 2352 34886 2408
rect 34942 2352 34947 2408
rect 30557 2350 34947 2352
rect 30557 2347 30623 2350
rect 34881 2347 34947 2350
rect 964 2240 75028 2264
rect 964 2176 1740 2240
rect 1804 2176 1820 2240
rect 1884 2236 1900 2240
rect 1964 2236 1980 2240
rect 2044 2236 2060 2240
rect 2124 2236 2140 2240
rect 1884 2176 1900 2180
rect 1964 2176 1980 2180
rect 2044 2176 2060 2180
rect 2124 2176 2140 2180
rect 2204 2176 2220 2240
rect 2284 2176 7740 2240
rect 7804 2176 7820 2240
rect 7884 2176 7900 2240
rect 7964 2176 7980 2240
rect 8044 2176 8060 2240
rect 8124 2176 8140 2240
rect 8204 2176 8220 2240
rect 8284 2236 13740 2240
rect 8284 2180 11864 2236
rect 11920 2180 11944 2236
rect 12000 2180 12024 2236
rect 12080 2180 12104 2236
rect 12160 2180 13740 2236
rect 8284 2176 13740 2180
rect 13804 2176 13820 2240
rect 13884 2176 13900 2240
rect 13964 2176 13980 2240
rect 14044 2176 14060 2240
rect 14124 2176 14140 2240
rect 14204 2176 14220 2240
rect 14284 2176 19740 2240
rect 19804 2176 19820 2240
rect 19884 2176 19900 2240
rect 19964 2176 19980 2240
rect 20044 2176 20060 2240
rect 20124 2176 20140 2240
rect 20204 2176 20220 2240
rect 20284 2236 25740 2240
rect 20284 2180 21864 2236
rect 21920 2180 21944 2236
rect 22000 2180 22024 2236
rect 22080 2180 22104 2236
rect 22160 2180 25740 2236
rect 20284 2176 25740 2180
rect 25804 2176 25820 2240
rect 25884 2176 25900 2240
rect 25964 2176 25980 2240
rect 26044 2176 26060 2240
rect 26124 2176 26140 2240
rect 26204 2176 26220 2240
rect 26284 2176 31740 2240
rect 31804 2176 31820 2240
rect 31884 2236 31900 2240
rect 31964 2236 31980 2240
rect 32044 2236 32060 2240
rect 32124 2236 32140 2240
rect 31884 2176 31900 2180
rect 31964 2176 31980 2180
rect 32044 2176 32060 2180
rect 32124 2176 32140 2180
rect 32204 2176 32220 2240
rect 32284 2176 37740 2240
rect 37804 2176 37820 2240
rect 37884 2176 37900 2240
rect 37964 2176 37980 2240
rect 38044 2176 38060 2240
rect 38124 2176 38140 2240
rect 38204 2176 38220 2240
rect 38284 2236 43740 2240
rect 38284 2180 41864 2236
rect 41920 2180 41944 2236
rect 42000 2180 42024 2236
rect 42080 2180 42104 2236
rect 42160 2180 43740 2236
rect 38284 2176 43740 2180
rect 43804 2176 43820 2240
rect 43884 2176 43900 2240
rect 43964 2176 43980 2240
rect 44044 2176 44060 2240
rect 44124 2176 44140 2240
rect 44204 2176 44220 2240
rect 44284 2176 49740 2240
rect 49804 2176 49820 2240
rect 49884 2176 49900 2240
rect 49964 2176 49980 2240
rect 50044 2176 50060 2240
rect 50124 2176 50140 2240
rect 50204 2176 50220 2240
rect 50284 2236 55740 2240
rect 50284 2180 51864 2236
rect 51920 2180 51944 2236
rect 52000 2180 52024 2236
rect 52080 2180 52104 2236
rect 52160 2180 55740 2236
rect 50284 2176 55740 2180
rect 55804 2176 55820 2240
rect 55884 2176 55900 2240
rect 55964 2176 55980 2240
rect 56044 2176 56060 2240
rect 56124 2176 56140 2240
rect 56204 2176 56220 2240
rect 56284 2176 61740 2240
rect 61804 2176 61820 2240
rect 61884 2236 61900 2240
rect 61964 2236 61980 2240
rect 62044 2236 62060 2240
rect 62124 2236 62140 2240
rect 61884 2176 61900 2180
rect 61964 2176 61980 2180
rect 62044 2176 62060 2180
rect 62124 2176 62140 2180
rect 62204 2176 62220 2240
rect 62284 2176 67740 2240
rect 67804 2176 67820 2240
rect 67884 2176 67900 2240
rect 67964 2176 67980 2240
rect 68044 2176 68060 2240
rect 68124 2176 68140 2240
rect 68204 2176 68220 2240
rect 68284 2236 73740 2240
rect 68284 2180 71864 2236
rect 71920 2180 71944 2236
rect 72000 2180 72024 2236
rect 72080 2180 72104 2236
rect 72160 2180 73740 2236
rect 68284 2176 73740 2180
rect 73804 2176 73820 2240
rect 73884 2176 73900 2240
rect 73964 2176 73980 2240
rect 74044 2176 74060 2240
rect 74124 2176 74140 2240
rect 74204 2176 74220 2240
rect 74284 2176 75028 2240
rect 964 2160 75028 2176
rect 964 2096 1740 2160
rect 1804 2096 1820 2160
rect 1884 2156 1900 2160
rect 1964 2156 1980 2160
rect 2044 2156 2060 2160
rect 2124 2156 2140 2160
rect 1884 2096 1900 2100
rect 1964 2096 1980 2100
rect 2044 2096 2060 2100
rect 2124 2096 2140 2100
rect 2204 2096 2220 2160
rect 2284 2096 7740 2160
rect 7804 2096 7820 2160
rect 7884 2096 7900 2160
rect 7964 2096 7980 2160
rect 8044 2096 8060 2160
rect 8124 2096 8140 2160
rect 8204 2096 8220 2160
rect 8284 2156 13740 2160
rect 8284 2100 11864 2156
rect 11920 2100 11944 2156
rect 12000 2100 12024 2156
rect 12080 2100 12104 2156
rect 12160 2100 13740 2156
rect 8284 2096 13740 2100
rect 13804 2096 13820 2160
rect 13884 2096 13900 2160
rect 13964 2096 13980 2160
rect 14044 2096 14060 2160
rect 14124 2096 14140 2160
rect 14204 2096 14220 2160
rect 14284 2096 19740 2160
rect 19804 2096 19820 2160
rect 19884 2096 19900 2160
rect 19964 2096 19980 2160
rect 20044 2096 20060 2160
rect 20124 2096 20140 2160
rect 20204 2096 20220 2160
rect 20284 2156 25740 2160
rect 20284 2100 21864 2156
rect 21920 2100 21944 2156
rect 22000 2100 22024 2156
rect 22080 2100 22104 2156
rect 22160 2100 25740 2156
rect 20284 2096 25740 2100
rect 25804 2096 25820 2160
rect 25884 2096 25900 2160
rect 25964 2096 25980 2160
rect 26044 2096 26060 2160
rect 26124 2096 26140 2160
rect 26204 2096 26220 2160
rect 26284 2096 31740 2160
rect 31804 2096 31820 2160
rect 31884 2156 31900 2160
rect 31964 2156 31980 2160
rect 32044 2156 32060 2160
rect 32124 2156 32140 2160
rect 31884 2096 31900 2100
rect 31964 2096 31980 2100
rect 32044 2096 32060 2100
rect 32124 2096 32140 2100
rect 32204 2096 32220 2160
rect 32284 2096 37740 2160
rect 37804 2096 37820 2160
rect 37884 2096 37900 2160
rect 37964 2096 37980 2160
rect 38044 2096 38060 2160
rect 38124 2096 38140 2160
rect 38204 2096 38220 2160
rect 38284 2156 43740 2160
rect 38284 2100 41864 2156
rect 41920 2100 41944 2156
rect 42000 2100 42024 2156
rect 42080 2100 42104 2156
rect 42160 2100 43740 2156
rect 38284 2096 43740 2100
rect 43804 2096 43820 2160
rect 43884 2096 43900 2160
rect 43964 2096 43980 2160
rect 44044 2096 44060 2160
rect 44124 2096 44140 2160
rect 44204 2096 44220 2160
rect 44284 2096 49740 2160
rect 49804 2096 49820 2160
rect 49884 2096 49900 2160
rect 49964 2096 49980 2160
rect 50044 2096 50060 2160
rect 50124 2096 50140 2160
rect 50204 2096 50220 2160
rect 50284 2156 55740 2160
rect 50284 2100 51864 2156
rect 51920 2100 51944 2156
rect 52000 2100 52024 2156
rect 52080 2100 52104 2156
rect 52160 2100 55740 2156
rect 50284 2096 55740 2100
rect 55804 2096 55820 2160
rect 55884 2096 55900 2160
rect 55964 2096 55980 2160
rect 56044 2096 56060 2160
rect 56124 2096 56140 2160
rect 56204 2096 56220 2160
rect 56284 2096 61740 2160
rect 61804 2096 61820 2160
rect 61884 2156 61900 2160
rect 61964 2156 61980 2160
rect 62044 2156 62060 2160
rect 62124 2156 62140 2160
rect 61884 2096 61900 2100
rect 61964 2096 61980 2100
rect 62044 2096 62060 2100
rect 62124 2096 62140 2100
rect 62204 2096 62220 2160
rect 62284 2096 67740 2160
rect 67804 2096 67820 2160
rect 67884 2096 67900 2160
rect 67964 2096 67980 2160
rect 68044 2096 68060 2160
rect 68124 2096 68140 2160
rect 68204 2096 68220 2160
rect 68284 2156 73740 2160
rect 68284 2100 71864 2156
rect 71920 2100 71944 2156
rect 72000 2100 72024 2156
rect 72080 2100 72104 2156
rect 72160 2100 73740 2156
rect 68284 2096 73740 2100
rect 73804 2096 73820 2160
rect 73884 2096 73900 2160
rect 73964 2096 73980 2160
rect 74044 2096 74060 2160
rect 74124 2096 74140 2160
rect 74204 2096 74220 2160
rect 74284 2096 75028 2160
rect 964 2080 75028 2096
rect 964 2016 1740 2080
rect 1804 2016 1820 2080
rect 1884 2076 1900 2080
rect 1964 2076 1980 2080
rect 2044 2076 2060 2080
rect 2124 2076 2140 2080
rect 1884 2016 1900 2020
rect 1964 2016 1980 2020
rect 2044 2016 2060 2020
rect 2124 2016 2140 2020
rect 2204 2016 2220 2080
rect 2284 2016 7740 2080
rect 7804 2016 7820 2080
rect 7884 2016 7900 2080
rect 7964 2016 7980 2080
rect 8044 2016 8060 2080
rect 8124 2016 8140 2080
rect 8204 2016 8220 2080
rect 8284 2076 13740 2080
rect 8284 2020 11864 2076
rect 11920 2020 11944 2076
rect 12000 2020 12024 2076
rect 12080 2020 12104 2076
rect 12160 2020 13740 2076
rect 8284 2016 13740 2020
rect 13804 2016 13820 2080
rect 13884 2016 13900 2080
rect 13964 2016 13980 2080
rect 14044 2016 14060 2080
rect 14124 2016 14140 2080
rect 14204 2016 14220 2080
rect 14284 2016 19740 2080
rect 19804 2016 19820 2080
rect 19884 2016 19900 2080
rect 19964 2016 19980 2080
rect 20044 2016 20060 2080
rect 20124 2016 20140 2080
rect 20204 2016 20220 2080
rect 20284 2076 25740 2080
rect 20284 2020 21864 2076
rect 21920 2020 21944 2076
rect 22000 2020 22024 2076
rect 22080 2020 22104 2076
rect 22160 2020 25740 2076
rect 20284 2016 25740 2020
rect 25804 2016 25820 2080
rect 25884 2016 25900 2080
rect 25964 2016 25980 2080
rect 26044 2016 26060 2080
rect 26124 2016 26140 2080
rect 26204 2016 26220 2080
rect 26284 2016 31740 2080
rect 31804 2016 31820 2080
rect 31884 2076 31900 2080
rect 31964 2076 31980 2080
rect 32044 2076 32060 2080
rect 32124 2076 32140 2080
rect 31884 2016 31900 2020
rect 31964 2016 31980 2020
rect 32044 2016 32060 2020
rect 32124 2016 32140 2020
rect 32204 2016 32220 2080
rect 32284 2016 37740 2080
rect 37804 2016 37820 2080
rect 37884 2016 37900 2080
rect 37964 2016 37980 2080
rect 38044 2016 38060 2080
rect 38124 2016 38140 2080
rect 38204 2016 38220 2080
rect 38284 2076 43740 2080
rect 38284 2020 41864 2076
rect 41920 2020 41944 2076
rect 42000 2020 42024 2076
rect 42080 2020 42104 2076
rect 42160 2020 43740 2076
rect 38284 2016 43740 2020
rect 43804 2016 43820 2080
rect 43884 2016 43900 2080
rect 43964 2016 43980 2080
rect 44044 2016 44060 2080
rect 44124 2016 44140 2080
rect 44204 2016 44220 2080
rect 44284 2016 49740 2080
rect 49804 2016 49820 2080
rect 49884 2016 49900 2080
rect 49964 2016 49980 2080
rect 50044 2016 50060 2080
rect 50124 2016 50140 2080
rect 50204 2016 50220 2080
rect 50284 2076 55740 2080
rect 50284 2020 51864 2076
rect 51920 2020 51944 2076
rect 52000 2020 52024 2076
rect 52080 2020 52104 2076
rect 52160 2020 55740 2076
rect 50284 2016 55740 2020
rect 55804 2016 55820 2080
rect 55884 2016 55900 2080
rect 55964 2016 55980 2080
rect 56044 2016 56060 2080
rect 56124 2016 56140 2080
rect 56204 2016 56220 2080
rect 56284 2016 61740 2080
rect 61804 2016 61820 2080
rect 61884 2076 61900 2080
rect 61964 2076 61980 2080
rect 62044 2076 62060 2080
rect 62124 2076 62140 2080
rect 61884 2016 61900 2020
rect 61964 2016 61980 2020
rect 62044 2016 62060 2020
rect 62124 2016 62140 2020
rect 62204 2016 62220 2080
rect 62284 2016 67740 2080
rect 67804 2016 67820 2080
rect 67884 2016 67900 2080
rect 67964 2016 67980 2080
rect 68044 2016 68060 2080
rect 68124 2016 68140 2080
rect 68204 2016 68220 2080
rect 68284 2076 73740 2080
rect 68284 2020 71864 2076
rect 71920 2020 71944 2076
rect 72000 2020 72024 2076
rect 72080 2020 72104 2076
rect 72160 2020 73740 2076
rect 68284 2016 73740 2020
rect 73804 2016 73820 2080
rect 73884 2016 73900 2080
rect 73964 2016 73980 2080
rect 74044 2016 74060 2080
rect 74124 2016 74140 2080
rect 74204 2016 74220 2080
rect 74284 2016 75028 2080
rect 964 2000 75028 2016
rect 964 1936 1740 2000
rect 1804 1936 1820 2000
rect 1884 1996 1900 2000
rect 1964 1996 1980 2000
rect 2044 1996 2060 2000
rect 2124 1996 2140 2000
rect 1884 1936 1900 1940
rect 1964 1936 1980 1940
rect 2044 1936 2060 1940
rect 2124 1936 2140 1940
rect 2204 1936 2220 2000
rect 2284 1936 7740 2000
rect 7804 1936 7820 2000
rect 7884 1936 7900 2000
rect 7964 1936 7980 2000
rect 8044 1936 8060 2000
rect 8124 1936 8140 2000
rect 8204 1936 8220 2000
rect 8284 1996 13740 2000
rect 8284 1940 11864 1996
rect 11920 1940 11944 1996
rect 12000 1940 12024 1996
rect 12080 1940 12104 1996
rect 12160 1940 13740 1996
rect 8284 1936 13740 1940
rect 13804 1936 13820 2000
rect 13884 1936 13900 2000
rect 13964 1936 13980 2000
rect 14044 1936 14060 2000
rect 14124 1936 14140 2000
rect 14204 1936 14220 2000
rect 14284 1936 19740 2000
rect 19804 1936 19820 2000
rect 19884 1936 19900 2000
rect 19964 1936 19980 2000
rect 20044 1936 20060 2000
rect 20124 1936 20140 2000
rect 20204 1936 20220 2000
rect 20284 1996 25740 2000
rect 20284 1940 21864 1996
rect 21920 1940 21944 1996
rect 22000 1940 22024 1996
rect 22080 1940 22104 1996
rect 22160 1940 25740 1996
rect 20284 1936 25740 1940
rect 25804 1936 25820 2000
rect 25884 1936 25900 2000
rect 25964 1936 25980 2000
rect 26044 1936 26060 2000
rect 26124 1936 26140 2000
rect 26204 1936 26220 2000
rect 26284 1936 31740 2000
rect 31804 1936 31820 2000
rect 31884 1996 31900 2000
rect 31964 1996 31980 2000
rect 32044 1996 32060 2000
rect 32124 1996 32140 2000
rect 31884 1936 31900 1940
rect 31964 1936 31980 1940
rect 32044 1936 32060 1940
rect 32124 1936 32140 1940
rect 32204 1936 32220 2000
rect 32284 1936 37740 2000
rect 37804 1936 37820 2000
rect 37884 1936 37900 2000
rect 37964 1936 37980 2000
rect 38044 1936 38060 2000
rect 38124 1936 38140 2000
rect 38204 1936 38220 2000
rect 38284 1996 43740 2000
rect 38284 1940 41864 1996
rect 41920 1940 41944 1996
rect 42000 1940 42024 1996
rect 42080 1940 42104 1996
rect 42160 1940 43740 1996
rect 38284 1936 43740 1940
rect 43804 1936 43820 2000
rect 43884 1936 43900 2000
rect 43964 1936 43980 2000
rect 44044 1936 44060 2000
rect 44124 1936 44140 2000
rect 44204 1936 44220 2000
rect 44284 1936 49740 2000
rect 49804 1936 49820 2000
rect 49884 1936 49900 2000
rect 49964 1936 49980 2000
rect 50044 1936 50060 2000
rect 50124 1936 50140 2000
rect 50204 1936 50220 2000
rect 50284 1996 55740 2000
rect 50284 1940 51864 1996
rect 51920 1940 51944 1996
rect 52000 1940 52024 1996
rect 52080 1940 52104 1996
rect 52160 1940 55740 1996
rect 50284 1936 55740 1940
rect 55804 1936 55820 2000
rect 55884 1936 55900 2000
rect 55964 1936 55980 2000
rect 56044 1936 56060 2000
rect 56124 1936 56140 2000
rect 56204 1936 56220 2000
rect 56284 1936 61740 2000
rect 61804 1936 61820 2000
rect 61884 1996 61900 2000
rect 61964 1996 61980 2000
rect 62044 1996 62060 2000
rect 62124 1996 62140 2000
rect 61884 1936 61900 1940
rect 61964 1936 61980 1940
rect 62044 1936 62060 1940
rect 62124 1936 62140 1940
rect 62204 1936 62220 2000
rect 62284 1936 67740 2000
rect 67804 1936 67820 2000
rect 67884 1936 67900 2000
rect 67964 1936 67980 2000
rect 68044 1936 68060 2000
rect 68124 1936 68140 2000
rect 68204 1936 68220 2000
rect 68284 1996 73740 2000
rect 68284 1940 71864 1996
rect 71920 1940 71944 1996
rect 72000 1940 72024 1996
rect 72080 1940 72104 1996
rect 72160 1940 73740 1996
rect 68284 1936 73740 1940
rect 73804 1936 73820 2000
rect 73884 1936 73900 2000
rect 73964 1936 73980 2000
rect 74044 1936 74060 2000
rect 74124 1936 74140 2000
rect 74204 1936 74220 2000
rect 74284 1936 75028 2000
rect 964 1912 75028 1936
rect 41137 1730 41203 1733
rect 47945 1730 48011 1733
rect 41137 1728 48011 1730
rect 41137 1672 41142 1728
rect 41198 1672 47950 1728
rect 48006 1672 48011 1728
rect 41137 1670 48011 1672
rect 41137 1667 41203 1670
rect 47945 1667 48011 1670
rect 33961 1322 34027 1325
rect 65558 1322 65564 1324
rect 33961 1320 65564 1322
rect 33961 1264 33966 1320
rect 34022 1264 65564 1320
rect 33961 1262 65564 1264
rect 33961 1259 34027 1262
rect 65558 1260 65564 1262
rect 65628 1260 65634 1324
<< via3 >>
rect 4740 84528 4804 84592
rect 4820 84528 4884 84592
rect 4900 84528 4964 84592
rect 4980 84528 5044 84592
rect 5060 84528 5124 84592
rect 5140 84528 5204 84592
rect 5220 84528 5284 84592
rect 10740 84528 10804 84592
rect 10820 84528 10884 84592
rect 10900 84528 10964 84592
rect 10980 84528 11044 84592
rect 11060 84528 11124 84592
rect 11140 84528 11204 84592
rect 11220 84528 11284 84592
rect 16740 84528 16804 84592
rect 16820 84528 16884 84592
rect 16900 84528 16964 84592
rect 16980 84528 17044 84592
rect 17060 84528 17124 84592
rect 17140 84588 17204 84592
rect 17220 84588 17284 84592
rect 17140 84532 17192 84588
rect 17192 84532 17204 84588
rect 17220 84532 17248 84588
rect 17248 84532 17284 84588
rect 17140 84528 17204 84532
rect 17220 84528 17284 84532
rect 22740 84528 22804 84592
rect 22820 84528 22884 84592
rect 22900 84528 22964 84592
rect 22980 84588 23044 84592
rect 22980 84532 23028 84588
rect 23028 84532 23044 84588
rect 22980 84528 23044 84532
rect 23060 84528 23124 84592
rect 23140 84528 23204 84592
rect 23220 84528 23284 84592
rect 28740 84588 28804 84592
rect 28740 84532 28752 84588
rect 28752 84532 28804 84588
rect 28740 84528 28804 84532
rect 28820 84528 28884 84592
rect 28900 84528 28964 84592
rect 28980 84528 29044 84592
rect 29060 84528 29124 84592
rect 29140 84528 29204 84592
rect 29220 84528 29284 84592
rect 34740 84528 34804 84592
rect 34820 84528 34884 84592
rect 34900 84528 34964 84592
rect 34980 84528 35044 84592
rect 35060 84528 35124 84592
rect 35140 84528 35204 84592
rect 35220 84528 35284 84592
rect 40740 84528 40804 84592
rect 40820 84528 40884 84592
rect 40900 84528 40964 84592
rect 40980 84528 41044 84592
rect 41060 84528 41124 84592
rect 41140 84528 41204 84592
rect 41220 84528 41284 84592
rect 46740 84528 46804 84592
rect 46820 84528 46884 84592
rect 46900 84528 46964 84592
rect 46980 84528 47044 84592
rect 47060 84528 47124 84592
rect 47140 84528 47204 84592
rect 47220 84528 47284 84592
rect 52740 84528 52804 84592
rect 52820 84528 52884 84592
rect 52900 84528 52964 84592
rect 52980 84528 53044 84592
rect 53060 84528 53124 84592
rect 53140 84528 53204 84592
rect 53220 84528 53284 84592
rect 58740 84528 58804 84592
rect 58820 84528 58884 84592
rect 58900 84528 58964 84592
rect 58980 84528 59044 84592
rect 59060 84528 59124 84592
rect 59140 84588 59204 84592
rect 59140 84532 59196 84588
rect 59196 84532 59204 84588
rect 59140 84528 59204 84532
rect 59220 84528 59284 84592
rect 64740 84528 64804 84592
rect 64820 84528 64884 84592
rect 64900 84528 64964 84592
rect 64980 84528 65044 84592
rect 65060 84528 65124 84592
rect 65140 84528 65204 84592
rect 65220 84528 65284 84592
rect 70740 84528 70804 84592
rect 70820 84528 70884 84592
rect 70900 84528 70964 84592
rect 70980 84528 71044 84592
rect 71060 84528 71124 84592
rect 71140 84528 71204 84592
rect 71220 84528 71284 84592
rect 4740 84448 4804 84512
rect 4820 84448 4884 84512
rect 4900 84448 4964 84512
rect 4980 84448 5044 84512
rect 5060 84448 5124 84512
rect 5140 84448 5204 84512
rect 5220 84448 5284 84512
rect 10740 84448 10804 84512
rect 10820 84448 10884 84512
rect 10900 84448 10964 84512
rect 10980 84448 11044 84512
rect 11060 84448 11124 84512
rect 11140 84448 11204 84512
rect 11220 84448 11284 84512
rect 16740 84448 16804 84512
rect 16820 84448 16884 84512
rect 16900 84448 16964 84512
rect 16980 84448 17044 84512
rect 17060 84448 17124 84512
rect 17140 84508 17204 84512
rect 17220 84508 17284 84512
rect 17140 84452 17192 84508
rect 17192 84452 17204 84508
rect 17220 84452 17248 84508
rect 17248 84452 17284 84508
rect 17140 84448 17204 84452
rect 17220 84448 17284 84452
rect 22740 84448 22804 84512
rect 22820 84448 22884 84512
rect 22900 84448 22964 84512
rect 22980 84508 23044 84512
rect 22980 84452 23028 84508
rect 23028 84452 23044 84508
rect 22980 84448 23044 84452
rect 23060 84448 23124 84512
rect 23140 84448 23204 84512
rect 23220 84448 23284 84512
rect 28740 84508 28804 84512
rect 28740 84452 28752 84508
rect 28752 84452 28804 84508
rect 28740 84448 28804 84452
rect 28820 84448 28884 84512
rect 28900 84448 28964 84512
rect 28980 84448 29044 84512
rect 29060 84448 29124 84512
rect 29140 84448 29204 84512
rect 29220 84448 29284 84512
rect 34740 84448 34804 84512
rect 34820 84448 34884 84512
rect 34900 84448 34964 84512
rect 34980 84448 35044 84512
rect 35060 84448 35124 84512
rect 35140 84448 35204 84512
rect 35220 84448 35284 84512
rect 40740 84448 40804 84512
rect 40820 84448 40884 84512
rect 40900 84448 40964 84512
rect 40980 84448 41044 84512
rect 41060 84448 41124 84512
rect 41140 84448 41204 84512
rect 41220 84448 41284 84512
rect 46740 84448 46804 84512
rect 46820 84448 46884 84512
rect 46900 84448 46964 84512
rect 46980 84448 47044 84512
rect 47060 84448 47124 84512
rect 47140 84448 47204 84512
rect 47220 84448 47284 84512
rect 52740 84448 52804 84512
rect 52820 84448 52884 84512
rect 52900 84448 52964 84512
rect 52980 84448 53044 84512
rect 53060 84448 53124 84512
rect 53140 84448 53204 84512
rect 53220 84448 53284 84512
rect 58740 84448 58804 84512
rect 58820 84448 58884 84512
rect 58900 84448 58964 84512
rect 58980 84448 59044 84512
rect 59060 84448 59124 84512
rect 59140 84508 59204 84512
rect 59140 84452 59196 84508
rect 59196 84452 59204 84508
rect 59140 84448 59204 84452
rect 59220 84448 59284 84512
rect 64740 84448 64804 84512
rect 64820 84448 64884 84512
rect 64900 84448 64964 84512
rect 64980 84448 65044 84512
rect 65060 84448 65124 84512
rect 65140 84448 65204 84512
rect 65220 84448 65284 84512
rect 70740 84448 70804 84512
rect 70820 84448 70884 84512
rect 70900 84448 70964 84512
rect 70980 84448 71044 84512
rect 71060 84448 71124 84512
rect 71140 84448 71204 84512
rect 71220 84448 71284 84512
rect 4740 84368 4804 84432
rect 4820 84368 4884 84432
rect 4900 84368 4964 84432
rect 4980 84368 5044 84432
rect 5060 84368 5124 84432
rect 5140 84368 5204 84432
rect 5220 84368 5284 84432
rect 10740 84368 10804 84432
rect 10820 84368 10884 84432
rect 10900 84368 10964 84432
rect 10980 84368 11044 84432
rect 11060 84368 11124 84432
rect 11140 84368 11204 84432
rect 11220 84368 11284 84432
rect 16740 84368 16804 84432
rect 16820 84368 16884 84432
rect 16900 84368 16964 84432
rect 16980 84368 17044 84432
rect 17060 84368 17124 84432
rect 17140 84428 17204 84432
rect 17220 84428 17284 84432
rect 17140 84372 17192 84428
rect 17192 84372 17204 84428
rect 17220 84372 17248 84428
rect 17248 84372 17284 84428
rect 17140 84368 17204 84372
rect 17220 84368 17284 84372
rect 22740 84368 22804 84432
rect 22820 84368 22884 84432
rect 22900 84368 22964 84432
rect 22980 84428 23044 84432
rect 22980 84372 23028 84428
rect 23028 84372 23044 84428
rect 22980 84368 23044 84372
rect 23060 84368 23124 84432
rect 23140 84368 23204 84432
rect 23220 84368 23284 84432
rect 28740 84428 28804 84432
rect 28740 84372 28752 84428
rect 28752 84372 28804 84428
rect 28740 84368 28804 84372
rect 28820 84368 28884 84432
rect 28900 84368 28964 84432
rect 28980 84368 29044 84432
rect 29060 84368 29124 84432
rect 29140 84368 29204 84432
rect 29220 84368 29284 84432
rect 34740 84368 34804 84432
rect 34820 84368 34884 84432
rect 34900 84368 34964 84432
rect 34980 84368 35044 84432
rect 35060 84368 35124 84432
rect 35140 84368 35204 84432
rect 35220 84368 35284 84432
rect 40740 84368 40804 84432
rect 40820 84368 40884 84432
rect 40900 84368 40964 84432
rect 40980 84368 41044 84432
rect 41060 84368 41124 84432
rect 41140 84368 41204 84432
rect 41220 84368 41284 84432
rect 46740 84368 46804 84432
rect 46820 84368 46884 84432
rect 46900 84368 46964 84432
rect 46980 84368 47044 84432
rect 47060 84368 47124 84432
rect 47140 84368 47204 84432
rect 47220 84368 47284 84432
rect 52740 84368 52804 84432
rect 52820 84368 52884 84432
rect 52900 84368 52964 84432
rect 52980 84368 53044 84432
rect 53060 84368 53124 84432
rect 53140 84368 53204 84432
rect 53220 84368 53284 84432
rect 58740 84368 58804 84432
rect 58820 84368 58884 84432
rect 58900 84368 58964 84432
rect 58980 84368 59044 84432
rect 59060 84368 59124 84432
rect 59140 84428 59204 84432
rect 59140 84372 59196 84428
rect 59196 84372 59204 84428
rect 59140 84368 59204 84372
rect 59220 84368 59284 84432
rect 64740 84368 64804 84432
rect 64820 84368 64884 84432
rect 64900 84368 64964 84432
rect 64980 84368 65044 84432
rect 65060 84368 65124 84432
rect 65140 84368 65204 84432
rect 65220 84368 65284 84432
rect 70740 84368 70804 84432
rect 70820 84368 70884 84432
rect 70900 84368 70964 84432
rect 70980 84368 71044 84432
rect 71060 84368 71124 84432
rect 71140 84368 71204 84432
rect 71220 84368 71284 84432
rect 4740 84288 4804 84352
rect 4820 84288 4884 84352
rect 4900 84288 4964 84352
rect 4980 84288 5044 84352
rect 5060 84288 5124 84352
rect 5140 84288 5204 84352
rect 5220 84288 5284 84352
rect 10740 84288 10804 84352
rect 10820 84288 10884 84352
rect 10900 84288 10964 84352
rect 10980 84288 11044 84352
rect 11060 84288 11124 84352
rect 11140 84288 11204 84352
rect 11220 84288 11284 84352
rect 16740 84288 16804 84352
rect 16820 84288 16884 84352
rect 16900 84288 16964 84352
rect 16980 84288 17044 84352
rect 17060 84288 17124 84352
rect 17140 84348 17204 84352
rect 17220 84348 17284 84352
rect 17140 84292 17192 84348
rect 17192 84292 17204 84348
rect 17220 84292 17248 84348
rect 17248 84292 17284 84348
rect 17140 84288 17204 84292
rect 17220 84288 17284 84292
rect 22740 84288 22804 84352
rect 22820 84288 22884 84352
rect 22900 84288 22964 84352
rect 22980 84348 23044 84352
rect 22980 84292 23028 84348
rect 23028 84292 23044 84348
rect 22980 84288 23044 84292
rect 23060 84288 23124 84352
rect 23140 84288 23204 84352
rect 23220 84288 23284 84352
rect 28740 84348 28804 84352
rect 28740 84292 28752 84348
rect 28752 84292 28804 84348
rect 28740 84288 28804 84292
rect 28820 84288 28884 84352
rect 28900 84288 28964 84352
rect 28980 84288 29044 84352
rect 29060 84288 29124 84352
rect 29140 84288 29204 84352
rect 29220 84288 29284 84352
rect 34740 84288 34804 84352
rect 34820 84288 34884 84352
rect 34900 84288 34964 84352
rect 34980 84288 35044 84352
rect 35060 84288 35124 84352
rect 35140 84288 35204 84352
rect 35220 84288 35284 84352
rect 40740 84288 40804 84352
rect 40820 84288 40884 84352
rect 40900 84288 40964 84352
rect 40980 84288 41044 84352
rect 41060 84288 41124 84352
rect 41140 84288 41204 84352
rect 41220 84288 41284 84352
rect 46740 84288 46804 84352
rect 46820 84288 46884 84352
rect 46900 84288 46964 84352
rect 46980 84288 47044 84352
rect 47060 84288 47124 84352
rect 47140 84288 47204 84352
rect 47220 84288 47284 84352
rect 52740 84288 52804 84352
rect 52820 84288 52884 84352
rect 52900 84288 52964 84352
rect 52980 84288 53044 84352
rect 53060 84288 53124 84352
rect 53140 84288 53204 84352
rect 53220 84288 53284 84352
rect 58740 84288 58804 84352
rect 58820 84288 58884 84352
rect 58900 84288 58964 84352
rect 58980 84288 59044 84352
rect 59060 84288 59124 84352
rect 59140 84348 59204 84352
rect 59140 84292 59196 84348
rect 59196 84292 59204 84348
rect 59140 84288 59204 84292
rect 59220 84288 59284 84352
rect 64740 84288 64804 84352
rect 64820 84288 64884 84352
rect 64900 84288 64964 84352
rect 64980 84288 65044 84352
rect 65060 84288 65124 84352
rect 65140 84288 65204 84352
rect 65220 84288 65284 84352
rect 70740 84288 70804 84352
rect 70820 84288 70884 84352
rect 70900 84288 70964 84352
rect 70980 84288 71044 84352
rect 71060 84288 71124 84352
rect 71140 84288 71204 84352
rect 71220 84288 71284 84352
rect 1740 82176 1804 82240
rect 1820 82176 1884 82240
rect 1900 82176 1964 82240
rect 1980 82176 2044 82240
rect 2060 82176 2124 82240
rect 2140 82176 2204 82240
rect 2220 82236 2284 82240
rect 2220 82180 2276 82236
rect 2276 82180 2284 82236
rect 2220 82176 2284 82180
rect 7740 82176 7804 82240
rect 7820 82176 7884 82240
rect 7900 82176 7964 82240
rect 7980 82176 8044 82240
rect 8060 82176 8124 82240
rect 8140 82176 8204 82240
rect 8220 82176 8284 82240
rect 13740 82176 13804 82240
rect 13820 82176 13884 82240
rect 13900 82176 13964 82240
rect 13980 82176 14044 82240
rect 14060 82176 14124 82240
rect 14140 82236 14204 82240
rect 14140 82180 14155 82236
rect 14155 82180 14204 82236
rect 14140 82176 14204 82180
rect 14220 82176 14284 82240
rect 19740 82176 19804 82240
rect 19820 82176 19884 82240
rect 19900 82236 19964 82240
rect 19980 82236 20044 82240
rect 19900 82180 19935 82236
rect 19935 82180 19964 82236
rect 19980 82180 19991 82236
rect 19991 82180 20044 82236
rect 19900 82176 19964 82180
rect 19980 82176 20044 82180
rect 20060 82176 20124 82240
rect 20140 82176 20204 82240
rect 20220 82176 20284 82240
rect 25740 82236 25804 82240
rect 25740 82180 25771 82236
rect 25771 82180 25804 82236
rect 25740 82176 25804 82180
rect 25820 82176 25884 82240
rect 25900 82176 25964 82240
rect 25980 82176 26044 82240
rect 26060 82176 26124 82240
rect 26140 82176 26204 82240
rect 26220 82176 26284 82240
rect 31740 82176 31804 82240
rect 31820 82176 31884 82240
rect 31900 82176 31964 82240
rect 31980 82176 32044 82240
rect 32060 82176 32124 82240
rect 32140 82176 32204 82240
rect 32220 82176 32284 82240
rect 37740 82176 37804 82240
rect 37820 82176 37884 82240
rect 37900 82176 37964 82240
rect 37980 82176 38044 82240
rect 38060 82176 38124 82240
rect 38140 82176 38204 82240
rect 38220 82176 38284 82240
rect 43740 82176 43804 82240
rect 43820 82176 43884 82240
rect 43900 82176 43964 82240
rect 43980 82176 44044 82240
rect 44060 82176 44124 82240
rect 44140 82176 44204 82240
rect 44220 82176 44284 82240
rect 49740 82236 49804 82240
rect 49820 82236 49884 82240
rect 49740 82180 49754 82236
rect 49754 82180 49804 82236
rect 49820 82180 49834 82236
rect 49834 82180 49884 82236
rect 49740 82176 49804 82180
rect 49820 82176 49884 82180
rect 49900 82176 49964 82240
rect 49980 82176 50044 82240
rect 50060 82176 50124 82240
rect 50140 82176 50204 82240
rect 50220 82176 50284 82240
rect 55740 82176 55804 82240
rect 55820 82176 55884 82240
rect 55900 82176 55964 82240
rect 55980 82176 56044 82240
rect 56060 82176 56124 82240
rect 56140 82176 56204 82240
rect 56220 82176 56284 82240
rect 61740 82176 61804 82240
rect 61820 82176 61884 82240
rect 61900 82176 61964 82240
rect 61980 82176 62044 82240
rect 62060 82176 62124 82240
rect 62140 82176 62204 82240
rect 62220 82176 62284 82240
rect 67740 82176 67804 82240
rect 67820 82176 67884 82240
rect 67900 82176 67964 82240
rect 67980 82176 68044 82240
rect 68060 82176 68124 82240
rect 68140 82176 68204 82240
rect 68220 82176 68284 82240
rect 73740 82176 73804 82240
rect 73820 82176 73884 82240
rect 73900 82176 73964 82240
rect 73980 82176 74044 82240
rect 74060 82176 74124 82240
rect 74140 82176 74204 82240
rect 74220 82176 74284 82240
rect 1740 82096 1804 82160
rect 1820 82096 1884 82160
rect 1900 82096 1964 82160
rect 1980 82096 2044 82160
rect 2060 82096 2124 82160
rect 2140 82096 2204 82160
rect 2220 82156 2284 82160
rect 2220 82100 2276 82156
rect 2276 82100 2284 82156
rect 2220 82096 2284 82100
rect 7740 82096 7804 82160
rect 7820 82096 7884 82160
rect 7900 82096 7964 82160
rect 7980 82096 8044 82160
rect 8060 82096 8124 82160
rect 8140 82096 8204 82160
rect 8220 82096 8284 82160
rect 13740 82096 13804 82160
rect 13820 82096 13884 82160
rect 13900 82096 13964 82160
rect 13980 82096 14044 82160
rect 14060 82096 14124 82160
rect 14140 82156 14204 82160
rect 14140 82100 14155 82156
rect 14155 82100 14204 82156
rect 14140 82096 14204 82100
rect 14220 82096 14284 82160
rect 19740 82096 19804 82160
rect 19820 82096 19884 82160
rect 19900 82156 19964 82160
rect 19980 82156 20044 82160
rect 19900 82100 19935 82156
rect 19935 82100 19964 82156
rect 19980 82100 19991 82156
rect 19991 82100 20044 82156
rect 19900 82096 19964 82100
rect 19980 82096 20044 82100
rect 20060 82096 20124 82160
rect 20140 82096 20204 82160
rect 20220 82096 20284 82160
rect 25740 82156 25804 82160
rect 25740 82100 25771 82156
rect 25771 82100 25804 82156
rect 25740 82096 25804 82100
rect 25820 82096 25884 82160
rect 25900 82096 25964 82160
rect 25980 82096 26044 82160
rect 26060 82096 26124 82160
rect 26140 82096 26204 82160
rect 26220 82096 26284 82160
rect 31740 82096 31804 82160
rect 31820 82096 31884 82160
rect 31900 82096 31964 82160
rect 31980 82096 32044 82160
rect 32060 82096 32124 82160
rect 32140 82096 32204 82160
rect 32220 82096 32284 82160
rect 37740 82096 37804 82160
rect 37820 82096 37884 82160
rect 37900 82096 37964 82160
rect 37980 82096 38044 82160
rect 38060 82096 38124 82160
rect 38140 82096 38204 82160
rect 38220 82096 38284 82160
rect 43740 82096 43804 82160
rect 43820 82096 43884 82160
rect 43900 82096 43964 82160
rect 43980 82096 44044 82160
rect 44060 82096 44124 82160
rect 44140 82096 44204 82160
rect 44220 82096 44284 82160
rect 49740 82156 49804 82160
rect 49820 82156 49884 82160
rect 49740 82100 49754 82156
rect 49754 82100 49804 82156
rect 49820 82100 49834 82156
rect 49834 82100 49884 82156
rect 49740 82096 49804 82100
rect 49820 82096 49884 82100
rect 49900 82096 49964 82160
rect 49980 82096 50044 82160
rect 50060 82096 50124 82160
rect 50140 82096 50204 82160
rect 50220 82096 50284 82160
rect 55740 82096 55804 82160
rect 55820 82096 55884 82160
rect 55900 82096 55964 82160
rect 55980 82096 56044 82160
rect 56060 82096 56124 82160
rect 56140 82096 56204 82160
rect 56220 82096 56284 82160
rect 61740 82096 61804 82160
rect 61820 82096 61884 82160
rect 61900 82096 61964 82160
rect 61980 82096 62044 82160
rect 62060 82096 62124 82160
rect 62140 82096 62204 82160
rect 62220 82096 62284 82160
rect 67740 82096 67804 82160
rect 67820 82096 67884 82160
rect 67900 82096 67964 82160
rect 67980 82096 68044 82160
rect 68060 82096 68124 82160
rect 68140 82096 68204 82160
rect 68220 82096 68284 82160
rect 73740 82096 73804 82160
rect 73820 82096 73884 82160
rect 73900 82096 73964 82160
rect 73980 82096 74044 82160
rect 74060 82096 74124 82160
rect 74140 82096 74204 82160
rect 74220 82096 74284 82160
rect 1740 82016 1804 82080
rect 1820 82016 1884 82080
rect 1900 82016 1964 82080
rect 1980 82016 2044 82080
rect 2060 82016 2124 82080
rect 2140 82016 2204 82080
rect 2220 82076 2284 82080
rect 2220 82020 2276 82076
rect 2276 82020 2284 82076
rect 2220 82016 2284 82020
rect 7740 82016 7804 82080
rect 7820 82016 7884 82080
rect 7900 82016 7964 82080
rect 7980 82016 8044 82080
rect 8060 82016 8124 82080
rect 8140 82016 8204 82080
rect 8220 82016 8284 82080
rect 13740 82016 13804 82080
rect 13820 82016 13884 82080
rect 13900 82016 13964 82080
rect 13980 82016 14044 82080
rect 14060 82016 14124 82080
rect 14140 82076 14204 82080
rect 14140 82020 14155 82076
rect 14155 82020 14204 82076
rect 14140 82016 14204 82020
rect 14220 82016 14284 82080
rect 19740 82016 19804 82080
rect 19820 82016 19884 82080
rect 19900 82076 19964 82080
rect 19980 82076 20044 82080
rect 19900 82020 19935 82076
rect 19935 82020 19964 82076
rect 19980 82020 19991 82076
rect 19991 82020 20044 82076
rect 19900 82016 19964 82020
rect 19980 82016 20044 82020
rect 20060 82016 20124 82080
rect 20140 82016 20204 82080
rect 20220 82016 20284 82080
rect 25740 82076 25804 82080
rect 25740 82020 25771 82076
rect 25771 82020 25804 82076
rect 25740 82016 25804 82020
rect 25820 82016 25884 82080
rect 25900 82016 25964 82080
rect 25980 82016 26044 82080
rect 26060 82016 26124 82080
rect 26140 82016 26204 82080
rect 26220 82016 26284 82080
rect 31740 82016 31804 82080
rect 31820 82016 31884 82080
rect 31900 82016 31964 82080
rect 31980 82016 32044 82080
rect 32060 82016 32124 82080
rect 32140 82016 32204 82080
rect 32220 82016 32284 82080
rect 37740 82016 37804 82080
rect 37820 82016 37884 82080
rect 37900 82016 37964 82080
rect 37980 82016 38044 82080
rect 38060 82016 38124 82080
rect 38140 82016 38204 82080
rect 38220 82016 38284 82080
rect 43740 82016 43804 82080
rect 43820 82016 43884 82080
rect 43900 82016 43964 82080
rect 43980 82016 44044 82080
rect 44060 82016 44124 82080
rect 44140 82016 44204 82080
rect 44220 82016 44284 82080
rect 49740 82076 49804 82080
rect 49820 82076 49884 82080
rect 49740 82020 49754 82076
rect 49754 82020 49804 82076
rect 49820 82020 49834 82076
rect 49834 82020 49884 82076
rect 49740 82016 49804 82020
rect 49820 82016 49884 82020
rect 49900 82016 49964 82080
rect 49980 82016 50044 82080
rect 50060 82016 50124 82080
rect 50140 82016 50204 82080
rect 50220 82016 50284 82080
rect 55740 82016 55804 82080
rect 55820 82016 55884 82080
rect 55900 82016 55964 82080
rect 55980 82016 56044 82080
rect 56060 82016 56124 82080
rect 56140 82016 56204 82080
rect 56220 82016 56284 82080
rect 61740 82016 61804 82080
rect 61820 82016 61884 82080
rect 61900 82016 61964 82080
rect 61980 82016 62044 82080
rect 62060 82016 62124 82080
rect 62140 82016 62204 82080
rect 62220 82016 62284 82080
rect 67740 82016 67804 82080
rect 67820 82016 67884 82080
rect 67900 82016 67964 82080
rect 67980 82016 68044 82080
rect 68060 82016 68124 82080
rect 68140 82016 68204 82080
rect 68220 82016 68284 82080
rect 73740 82016 73804 82080
rect 73820 82016 73884 82080
rect 73900 82016 73964 82080
rect 73980 82016 74044 82080
rect 74060 82016 74124 82080
rect 74140 82016 74204 82080
rect 74220 82016 74284 82080
rect 1740 81936 1804 82000
rect 1820 81936 1884 82000
rect 1900 81936 1964 82000
rect 1980 81936 2044 82000
rect 2060 81936 2124 82000
rect 2140 81936 2204 82000
rect 2220 81996 2284 82000
rect 2220 81940 2276 81996
rect 2276 81940 2284 81996
rect 2220 81936 2284 81940
rect 7740 81936 7804 82000
rect 7820 81936 7884 82000
rect 7900 81936 7964 82000
rect 7980 81936 8044 82000
rect 8060 81936 8124 82000
rect 8140 81936 8204 82000
rect 8220 81936 8284 82000
rect 13740 81936 13804 82000
rect 13820 81936 13884 82000
rect 13900 81936 13964 82000
rect 13980 81936 14044 82000
rect 14060 81936 14124 82000
rect 14140 81996 14204 82000
rect 14140 81940 14155 81996
rect 14155 81940 14204 81996
rect 14140 81936 14204 81940
rect 14220 81936 14284 82000
rect 19740 81936 19804 82000
rect 19820 81936 19884 82000
rect 19900 81996 19964 82000
rect 19980 81996 20044 82000
rect 19900 81940 19935 81996
rect 19935 81940 19964 81996
rect 19980 81940 19991 81996
rect 19991 81940 20044 81996
rect 19900 81936 19964 81940
rect 19980 81936 20044 81940
rect 20060 81936 20124 82000
rect 20140 81936 20204 82000
rect 20220 81936 20284 82000
rect 25740 81996 25804 82000
rect 25740 81940 25771 81996
rect 25771 81940 25804 81996
rect 25740 81936 25804 81940
rect 25820 81936 25884 82000
rect 25900 81936 25964 82000
rect 25980 81936 26044 82000
rect 26060 81936 26124 82000
rect 26140 81936 26204 82000
rect 26220 81936 26284 82000
rect 31740 81936 31804 82000
rect 31820 81936 31884 82000
rect 31900 81936 31964 82000
rect 31980 81936 32044 82000
rect 32060 81936 32124 82000
rect 32140 81936 32204 82000
rect 32220 81936 32284 82000
rect 37740 81936 37804 82000
rect 37820 81936 37884 82000
rect 37900 81936 37964 82000
rect 37980 81936 38044 82000
rect 38060 81936 38124 82000
rect 38140 81936 38204 82000
rect 38220 81936 38284 82000
rect 43740 81936 43804 82000
rect 43820 81936 43884 82000
rect 43900 81936 43964 82000
rect 43980 81936 44044 82000
rect 44060 81936 44124 82000
rect 44140 81936 44204 82000
rect 44220 81936 44284 82000
rect 49740 81996 49804 82000
rect 49820 81996 49884 82000
rect 49740 81940 49754 81996
rect 49754 81940 49804 81996
rect 49820 81940 49834 81996
rect 49834 81940 49884 81996
rect 49740 81936 49804 81940
rect 49820 81936 49884 81940
rect 49900 81936 49964 82000
rect 49980 81936 50044 82000
rect 50060 81936 50124 82000
rect 50140 81936 50204 82000
rect 50220 81936 50284 82000
rect 55740 81936 55804 82000
rect 55820 81936 55884 82000
rect 55900 81936 55964 82000
rect 55980 81936 56044 82000
rect 56060 81936 56124 82000
rect 56140 81936 56204 82000
rect 56220 81936 56284 82000
rect 61740 81936 61804 82000
rect 61820 81936 61884 82000
rect 61900 81936 61964 82000
rect 61980 81936 62044 82000
rect 62060 81936 62124 82000
rect 62140 81936 62204 82000
rect 62220 81936 62284 82000
rect 67740 81936 67804 82000
rect 67820 81936 67884 82000
rect 67900 81936 67964 82000
rect 67980 81936 68044 82000
rect 68060 81936 68124 82000
rect 68140 81936 68204 82000
rect 68220 81936 68284 82000
rect 73740 81936 73804 82000
rect 73820 81936 73884 82000
rect 73900 81936 73964 82000
rect 73980 81936 74044 82000
rect 74060 81936 74124 82000
rect 74140 81936 74204 82000
rect 74220 81936 74284 82000
rect 4740 74528 4804 74592
rect 4820 74528 4884 74592
rect 4900 74528 4964 74592
rect 4980 74528 5044 74592
rect 5060 74528 5124 74592
rect 5140 74528 5204 74592
rect 5220 74528 5284 74592
rect 10740 74528 10804 74592
rect 10820 74528 10884 74592
rect 10900 74528 10964 74592
rect 10980 74528 11044 74592
rect 11060 74528 11124 74592
rect 11140 74528 11204 74592
rect 11220 74528 11284 74592
rect 16740 74528 16804 74592
rect 16820 74528 16884 74592
rect 16900 74528 16964 74592
rect 16980 74528 17044 74592
rect 17060 74528 17124 74592
rect 17140 74588 17204 74592
rect 17220 74588 17284 74592
rect 17140 74532 17192 74588
rect 17192 74532 17204 74588
rect 17220 74532 17248 74588
rect 17248 74532 17284 74588
rect 17140 74528 17204 74532
rect 17220 74528 17284 74532
rect 22740 74528 22804 74592
rect 22820 74528 22884 74592
rect 22900 74528 22964 74592
rect 22980 74588 23044 74592
rect 22980 74532 23028 74588
rect 23028 74532 23044 74588
rect 22980 74528 23044 74532
rect 23060 74528 23124 74592
rect 23140 74528 23204 74592
rect 23220 74528 23284 74592
rect 28740 74588 28804 74592
rect 28740 74532 28752 74588
rect 28752 74532 28804 74588
rect 28740 74528 28804 74532
rect 28820 74528 28884 74592
rect 28900 74528 28964 74592
rect 28980 74528 29044 74592
rect 29060 74528 29124 74592
rect 29140 74528 29204 74592
rect 29220 74528 29284 74592
rect 34740 74528 34804 74592
rect 34820 74528 34884 74592
rect 34900 74528 34964 74592
rect 34980 74528 35044 74592
rect 35060 74528 35124 74592
rect 35140 74528 35204 74592
rect 35220 74528 35284 74592
rect 40740 74528 40804 74592
rect 40820 74528 40884 74592
rect 40900 74528 40964 74592
rect 40980 74528 41044 74592
rect 41060 74528 41124 74592
rect 41140 74528 41204 74592
rect 41220 74528 41284 74592
rect 46740 74528 46804 74592
rect 46820 74528 46884 74592
rect 46900 74528 46964 74592
rect 46980 74528 47044 74592
rect 47060 74528 47124 74592
rect 47140 74528 47204 74592
rect 47220 74528 47284 74592
rect 52740 74528 52804 74592
rect 52820 74528 52884 74592
rect 52900 74528 52964 74592
rect 52980 74528 53044 74592
rect 53060 74528 53124 74592
rect 53140 74528 53204 74592
rect 53220 74528 53284 74592
rect 58740 74528 58804 74592
rect 58820 74528 58884 74592
rect 58900 74528 58964 74592
rect 58980 74528 59044 74592
rect 59060 74528 59124 74592
rect 59140 74588 59204 74592
rect 59140 74532 59196 74588
rect 59196 74532 59204 74588
rect 59140 74528 59204 74532
rect 59220 74528 59284 74592
rect 64740 74528 64804 74592
rect 64820 74528 64884 74592
rect 64900 74528 64964 74592
rect 64980 74528 65044 74592
rect 65060 74528 65124 74592
rect 65140 74528 65204 74592
rect 65220 74528 65284 74592
rect 70740 74528 70804 74592
rect 70820 74528 70884 74592
rect 70900 74528 70964 74592
rect 70980 74528 71044 74592
rect 71060 74528 71124 74592
rect 71140 74528 71204 74592
rect 71220 74528 71284 74592
rect 4740 74448 4804 74512
rect 4820 74448 4884 74512
rect 4900 74448 4964 74512
rect 4980 74448 5044 74512
rect 5060 74448 5124 74512
rect 5140 74448 5204 74512
rect 5220 74448 5284 74512
rect 10740 74448 10804 74512
rect 10820 74448 10884 74512
rect 10900 74448 10964 74512
rect 10980 74448 11044 74512
rect 11060 74448 11124 74512
rect 11140 74448 11204 74512
rect 11220 74448 11284 74512
rect 16740 74448 16804 74512
rect 16820 74448 16884 74512
rect 16900 74448 16964 74512
rect 16980 74448 17044 74512
rect 17060 74448 17124 74512
rect 17140 74508 17204 74512
rect 17220 74508 17284 74512
rect 17140 74452 17192 74508
rect 17192 74452 17204 74508
rect 17220 74452 17248 74508
rect 17248 74452 17284 74508
rect 17140 74448 17204 74452
rect 17220 74448 17284 74452
rect 22740 74448 22804 74512
rect 22820 74448 22884 74512
rect 22900 74448 22964 74512
rect 22980 74508 23044 74512
rect 22980 74452 23028 74508
rect 23028 74452 23044 74508
rect 22980 74448 23044 74452
rect 23060 74448 23124 74512
rect 23140 74448 23204 74512
rect 23220 74448 23284 74512
rect 28740 74508 28804 74512
rect 28740 74452 28752 74508
rect 28752 74452 28804 74508
rect 28740 74448 28804 74452
rect 28820 74448 28884 74512
rect 28900 74448 28964 74512
rect 28980 74448 29044 74512
rect 29060 74448 29124 74512
rect 29140 74448 29204 74512
rect 29220 74448 29284 74512
rect 34740 74448 34804 74512
rect 34820 74448 34884 74512
rect 34900 74448 34964 74512
rect 34980 74448 35044 74512
rect 35060 74448 35124 74512
rect 35140 74448 35204 74512
rect 35220 74448 35284 74512
rect 40740 74448 40804 74512
rect 40820 74448 40884 74512
rect 40900 74448 40964 74512
rect 40980 74448 41044 74512
rect 41060 74448 41124 74512
rect 41140 74448 41204 74512
rect 41220 74448 41284 74512
rect 46740 74448 46804 74512
rect 46820 74448 46884 74512
rect 46900 74448 46964 74512
rect 46980 74448 47044 74512
rect 47060 74448 47124 74512
rect 47140 74448 47204 74512
rect 47220 74448 47284 74512
rect 52740 74448 52804 74512
rect 52820 74448 52884 74512
rect 52900 74448 52964 74512
rect 52980 74448 53044 74512
rect 53060 74448 53124 74512
rect 53140 74448 53204 74512
rect 53220 74448 53284 74512
rect 58740 74448 58804 74512
rect 58820 74448 58884 74512
rect 58900 74448 58964 74512
rect 58980 74448 59044 74512
rect 59060 74448 59124 74512
rect 59140 74508 59204 74512
rect 59140 74452 59196 74508
rect 59196 74452 59204 74508
rect 59140 74448 59204 74452
rect 59220 74448 59284 74512
rect 64740 74448 64804 74512
rect 64820 74448 64884 74512
rect 64900 74448 64964 74512
rect 64980 74448 65044 74512
rect 65060 74448 65124 74512
rect 65140 74448 65204 74512
rect 65220 74448 65284 74512
rect 70740 74448 70804 74512
rect 70820 74448 70884 74512
rect 70900 74448 70964 74512
rect 70980 74448 71044 74512
rect 71060 74448 71124 74512
rect 71140 74448 71204 74512
rect 71220 74448 71284 74512
rect 4740 74368 4804 74432
rect 4820 74368 4884 74432
rect 4900 74368 4964 74432
rect 4980 74368 5044 74432
rect 5060 74368 5124 74432
rect 5140 74368 5204 74432
rect 5220 74368 5284 74432
rect 10740 74368 10804 74432
rect 10820 74368 10884 74432
rect 10900 74368 10964 74432
rect 10980 74368 11044 74432
rect 11060 74368 11124 74432
rect 11140 74368 11204 74432
rect 11220 74368 11284 74432
rect 16740 74368 16804 74432
rect 16820 74368 16884 74432
rect 16900 74368 16964 74432
rect 16980 74368 17044 74432
rect 17060 74368 17124 74432
rect 17140 74428 17204 74432
rect 17220 74428 17284 74432
rect 17140 74372 17192 74428
rect 17192 74372 17204 74428
rect 17220 74372 17248 74428
rect 17248 74372 17284 74428
rect 17140 74368 17204 74372
rect 17220 74368 17284 74372
rect 22740 74368 22804 74432
rect 22820 74368 22884 74432
rect 22900 74368 22964 74432
rect 22980 74428 23044 74432
rect 22980 74372 23028 74428
rect 23028 74372 23044 74428
rect 22980 74368 23044 74372
rect 23060 74368 23124 74432
rect 23140 74368 23204 74432
rect 23220 74368 23284 74432
rect 28740 74428 28804 74432
rect 28740 74372 28752 74428
rect 28752 74372 28804 74428
rect 28740 74368 28804 74372
rect 28820 74368 28884 74432
rect 28900 74368 28964 74432
rect 28980 74368 29044 74432
rect 29060 74368 29124 74432
rect 29140 74368 29204 74432
rect 29220 74368 29284 74432
rect 34740 74368 34804 74432
rect 34820 74368 34884 74432
rect 34900 74368 34964 74432
rect 34980 74368 35044 74432
rect 35060 74368 35124 74432
rect 35140 74368 35204 74432
rect 35220 74368 35284 74432
rect 40740 74368 40804 74432
rect 40820 74368 40884 74432
rect 40900 74368 40964 74432
rect 40980 74368 41044 74432
rect 41060 74368 41124 74432
rect 41140 74368 41204 74432
rect 41220 74368 41284 74432
rect 46740 74368 46804 74432
rect 46820 74368 46884 74432
rect 46900 74368 46964 74432
rect 46980 74368 47044 74432
rect 47060 74368 47124 74432
rect 47140 74368 47204 74432
rect 47220 74368 47284 74432
rect 52740 74368 52804 74432
rect 52820 74368 52884 74432
rect 52900 74368 52964 74432
rect 52980 74368 53044 74432
rect 53060 74368 53124 74432
rect 53140 74368 53204 74432
rect 53220 74368 53284 74432
rect 58740 74368 58804 74432
rect 58820 74368 58884 74432
rect 58900 74368 58964 74432
rect 58980 74368 59044 74432
rect 59060 74368 59124 74432
rect 59140 74428 59204 74432
rect 59140 74372 59196 74428
rect 59196 74372 59204 74428
rect 59140 74368 59204 74372
rect 59220 74368 59284 74432
rect 64740 74368 64804 74432
rect 64820 74368 64884 74432
rect 64900 74368 64964 74432
rect 64980 74368 65044 74432
rect 65060 74368 65124 74432
rect 65140 74368 65204 74432
rect 65220 74368 65284 74432
rect 70740 74368 70804 74432
rect 70820 74368 70884 74432
rect 70900 74368 70964 74432
rect 70980 74368 71044 74432
rect 71060 74368 71124 74432
rect 71140 74368 71204 74432
rect 71220 74368 71284 74432
rect 4740 74288 4804 74352
rect 4820 74288 4884 74352
rect 4900 74288 4964 74352
rect 4980 74288 5044 74352
rect 5060 74288 5124 74352
rect 5140 74288 5204 74352
rect 5220 74288 5284 74352
rect 10740 74288 10804 74352
rect 10820 74288 10884 74352
rect 10900 74288 10964 74352
rect 10980 74288 11044 74352
rect 11060 74288 11124 74352
rect 11140 74288 11204 74352
rect 11220 74288 11284 74352
rect 16740 74288 16804 74352
rect 16820 74288 16884 74352
rect 16900 74288 16964 74352
rect 16980 74288 17044 74352
rect 17060 74288 17124 74352
rect 17140 74348 17204 74352
rect 17220 74348 17284 74352
rect 17140 74292 17192 74348
rect 17192 74292 17204 74348
rect 17220 74292 17248 74348
rect 17248 74292 17284 74348
rect 17140 74288 17204 74292
rect 17220 74288 17284 74292
rect 22740 74288 22804 74352
rect 22820 74288 22884 74352
rect 22900 74288 22964 74352
rect 22980 74348 23044 74352
rect 22980 74292 23028 74348
rect 23028 74292 23044 74348
rect 22980 74288 23044 74292
rect 23060 74288 23124 74352
rect 23140 74288 23204 74352
rect 23220 74288 23284 74352
rect 28740 74348 28804 74352
rect 28740 74292 28752 74348
rect 28752 74292 28804 74348
rect 28740 74288 28804 74292
rect 28820 74288 28884 74352
rect 28900 74288 28964 74352
rect 28980 74288 29044 74352
rect 29060 74288 29124 74352
rect 29140 74288 29204 74352
rect 29220 74288 29284 74352
rect 34740 74288 34804 74352
rect 34820 74288 34884 74352
rect 34900 74288 34964 74352
rect 34980 74288 35044 74352
rect 35060 74288 35124 74352
rect 35140 74288 35204 74352
rect 35220 74288 35284 74352
rect 40740 74288 40804 74352
rect 40820 74288 40884 74352
rect 40900 74288 40964 74352
rect 40980 74288 41044 74352
rect 41060 74288 41124 74352
rect 41140 74288 41204 74352
rect 41220 74288 41284 74352
rect 46740 74288 46804 74352
rect 46820 74288 46884 74352
rect 46900 74288 46964 74352
rect 46980 74288 47044 74352
rect 47060 74288 47124 74352
rect 47140 74288 47204 74352
rect 47220 74288 47284 74352
rect 52740 74288 52804 74352
rect 52820 74288 52884 74352
rect 52900 74288 52964 74352
rect 52980 74288 53044 74352
rect 53060 74288 53124 74352
rect 53140 74288 53204 74352
rect 53220 74288 53284 74352
rect 58740 74288 58804 74352
rect 58820 74288 58884 74352
rect 58900 74288 58964 74352
rect 58980 74288 59044 74352
rect 59060 74288 59124 74352
rect 59140 74348 59204 74352
rect 59140 74292 59196 74348
rect 59196 74292 59204 74348
rect 59140 74288 59204 74292
rect 59220 74288 59284 74352
rect 64740 74288 64804 74352
rect 64820 74288 64884 74352
rect 64900 74288 64964 74352
rect 64980 74288 65044 74352
rect 65060 74288 65124 74352
rect 65140 74288 65204 74352
rect 65220 74288 65284 74352
rect 70740 74288 70804 74352
rect 70820 74288 70884 74352
rect 70900 74288 70964 74352
rect 70980 74288 71044 74352
rect 71060 74288 71124 74352
rect 71140 74288 71204 74352
rect 71220 74288 71284 74352
rect 1740 72176 1804 72240
rect 1820 72176 1884 72240
rect 1900 72176 1964 72240
rect 1980 72176 2044 72240
rect 2060 72176 2124 72240
rect 2140 72176 2204 72240
rect 2220 72236 2284 72240
rect 2220 72180 2276 72236
rect 2276 72180 2284 72236
rect 2220 72176 2284 72180
rect 7740 72176 7804 72240
rect 7820 72176 7884 72240
rect 7900 72176 7964 72240
rect 7980 72176 8044 72240
rect 8060 72176 8124 72240
rect 8140 72176 8204 72240
rect 8220 72176 8284 72240
rect 13740 72176 13804 72240
rect 13820 72176 13884 72240
rect 13900 72176 13964 72240
rect 13980 72176 14044 72240
rect 14060 72176 14124 72240
rect 14140 72236 14204 72240
rect 14140 72180 14155 72236
rect 14155 72180 14204 72236
rect 14140 72176 14204 72180
rect 14220 72176 14284 72240
rect 19740 72176 19804 72240
rect 19820 72176 19884 72240
rect 19900 72236 19964 72240
rect 19980 72236 20044 72240
rect 19900 72180 19935 72236
rect 19935 72180 19964 72236
rect 19980 72180 19991 72236
rect 19991 72180 20044 72236
rect 19900 72176 19964 72180
rect 19980 72176 20044 72180
rect 20060 72176 20124 72240
rect 20140 72176 20204 72240
rect 20220 72176 20284 72240
rect 25740 72236 25804 72240
rect 25740 72180 25771 72236
rect 25771 72180 25804 72236
rect 25740 72176 25804 72180
rect 25820 72176 25884 72240
rect 25900 72176 25964 72240
rect 25980 72176 26044 72240
rect 26060 72176 26124 72240
rect 26140 72176 26204 72240
rect 26220 72176 26284 72240
rect 31740 72176 31804 72240
rect 31820 72176 31884 72240
rect 31900 72176 31964 72240
rect 31980 72176 32044 72240
rect 32060 72176 32124 72240
rect 32140 72176 32204 72240
rect 32220 72176 32284 72240
rect 37740 72176 37804 72240
rect 37820 72176 37884 72240
rect 37900 72176 37964 72240
rect 37980 72176 38044 72240
rect 38060 72176 38124 72240
rect 38140 72176 38204 72240
rect 38220 72176 38284 72240
rect 43740 72176 43804 72240
rect 43820 72176 43884 72240
rect 43900 72176 43964 72240
rect 43980 72176 44044 72240
rect 44060 72176 44124 72240
rect 44140 72176 44204 72240
rect 44220 72176 44284 72240
rect 49740 72236 49804 72240
rect 49820 72236 49884 72240
rect 49740 72180 49754 72236
rect 49754 72180 49804 72236
rect 49820 72180 49834 72236
rect 49834 72180 49884 72236
rect 49740 72176 49804 72180
rect 49820 72176 49884 72180
rect 49900 72176 49964 72240
rect 49980 72176 50044 72240
rect 50060 72176 50124 72240
rect 50140 72176 50204 72240
rect 50220 72176 50284 72240
rect 55740 72176 55804 72240
rect 55820 72176 55884 72240
rect 55900 72176 55964 72240
rect 55980 72176 56044 72240
rect 56060 72176 56124 72240
rect 56140 72176 56204 72240
rect 56220 72176 56284 72240
rect 61740 72176 61804 72240
rect 61820 72176 61884 72240
rect 61900 72176 61964 72240
rect 61980 72176 62044 72240
rect 62060 72176 62124 72240
rect 62140 72176 62204 72240
rect 62220 72176 62284 72240
rect 67740 72176 67804 72240
rect 67820 72176 67884 72240
rect 67900 72176 67964 72240
rect 67980 72176 68044 72240
rect 68060 72176 68124 72240
rect 68140 72176 68204 72240
rect 68220 72176 68284 72240
rect 73740 72176 73804 72240
rect 73820 72176 73884 72240
rect 73900 72176 73964 72240
rect 73980 72176 74044 72240
rect 74060 72176 74124 72240
rect 74140 72176 74204 72240
rect 74220 72176 74284 72240
rect 1740 72096 1804 72160
rect 1820 72096 1884 72160
rect 1900 72096 1964 72160
rect 1980 72096 2044 72160
rect 2060 72096 2124 72160
rect 2140 72096 2204 72160
rect 2220 72156 2284 72160
rect 2220 72100 2276 72156
rect 2276 72100 2284 72156
rect 2220 72096 2284 72100
rect 7740 72096 7804 72160
rect 7820 72096 7884 72160
rect 7900 72096 7964 72160
rect 7980 72096 8044 72160
rect 8060 72096 8124 72160
rect 8140 72096 8204 72160
rect 8220 72096 8284 72160
rect 13740 72096 13804 72160
rect 13820 72096 13884 72160
rect 13900 72096 13964 72160
rect 13980 72096 14044 72160
rect 14060 72096 14124 72160
rect 14140 72156 14204 72160
rect 14140 72100 14155 72156
rect 14155 72100 14204 72156
rect 14140 72096 14204 72100
rect 14220 72096 14284 72160
rect 19740 72096 19804 72160
rect 19820 72096 19884 72160
rect 19900 72156 19964 72160
rect 19980 72156 20044 72160
rect 19900 72100 19935 72156
rect 19935 72100 19964 72156
rect 19980 72100 19991 72156
rect 19991 72100 20044 72156
rect 19900 72096 19964 72100
rect 19980 72096 20044 72100
rect 20060 72096 20124 72160
rect 20140 72096 20204 72160
rect 20220 72096 20284 72160
rect 25740 72156 25804 72160
rect 25740 72100 25771 72156
rect 25771 72100 25804 72156
rect 25740 72096 25804 72100
rect 25820 72096 25884 72160
rect 25900 72096 25964 72160
rect 25980 72096 26044 72160
rect 26060 72096 26124 72160
rect 26140 72096 26204 72160
rect 26220 72096 26284 72160
rect 31740 72096 31804 72160
rect 31820 72096 31884 72160
rect 31900 72096 31964 72160
rect 31980 72096 32044 72160
rect 32060 72096 32124 72160
rect 32140 72096 32204 72160
rect 32220 72096 32284 72160
rect 37740 72096 37804 72160
rect 37820 72096 37884 72160
rect 37900 72096 37964 72160
rect 37980 72096 38044 72160
rect 38060 72096 38124 72160
rect 38140 72096 38204 72160
rect 38220 72096 38284 72160
rect 43740 72096 43804 72160
rect 43820 72096 43884 72160
rect 43900 72096 43964 72160
rect 43980 72096 44044 72160
rect 44060 72096 44124 72160
rect 44140 72096 44204 72160
rect 44220 72096 44284 72160
rect 49740 72156 49804 72160
rect 49820 72156 49884 72160
rect 49740 72100 49754 72156
rect 49754 72100 49804 72156
rect 49820 72100 49834 72156
rect 49834 72100 49884 72156
rect 49740 72096 49804 72100
rect 49820 72096 49884 72100
rect 49900 72096 49964 72160
rect 49980 72096 50044 72160
rect 50060 72096 50124 72160
rect 50140 72096 50204 72160
rect 50220 72096 50284 72160
rect 55740 72096 55804 72160
rect 55820 72096 55884 72160
rect 55900 72096 55964 72160
rect 55980 72096 56044 72160
rect 56060 72096 56124 72160
rect 56140 72096 56204 72160
rect 56220 72096 56284 72160
rect 61740 72096 61804 72160
rect 61820 72096 61884 72160
rect 61900 72096 61964 72160
rect 61980 72096 62044 72160
rect 62060 72096 62124 72160
rect 62140 72096 62204 72160
rect 62220 72096 62284 72160
rect 67740 72096 67804 72160
rect 67820 72096 67884 72160
rect 67900 72096 67964 72160
rect 67980 72096 68044 72160
rect 68060 72096 68124 72160
rect 68140 72096 68204 72160
rect 68220 72096 68284 72160
rect 73740 72096 73804 72160
rect 73820 72096 73884 72160
rect 73900 72096 73964 72160
rect 73980 72096 74044 72160
rect 74060 72096 74124 72160
rect 74140 72096 74204 72160
rect 74220 72096 74284 72160
rect 1740 72016 1804 72080
rect 1820 72016 1884 72080
rect 1900 72016 1964 72080
rect 1980 72016 2044 72080
rect 2060 72016 2124 72080
rect 2140 72016 2204 72080
rect 2220 72076 2284 72080
rect 2220 72020 2276 72076
rect 2276 72020 2284 72076
rect 2220 72016 2284 72020
rect 7740 72016 7804 72080
rect 7820 72016 7884 72080
rect 7900 72016 7964 72080
rect 7980 72016 8044 72080
rect 8060 72016 8124 72080
rect 8140 72016 8204 72080
rect 8220 72016 8284 72080
rect 13740 72016 13804 72080
rect 13820 72016 13884 72080
rect 13900 72016 13964 72080
rect 13980 72016 14044 72080
rect 14060 72016 14124 72080
rect 14140 72076 14204 72080
rect 14140 72020 14155 72076
rect 14155 72020 14204 72076
rect 14140 72016 14204 72020
rect 14220 72016 14284 72080
rect 19740 72016 19804 72080
rect 19820 72016 19884 72080
rect 19900 72076 19964 72080
rect 19980 72076 20044 72080
rect 19900 72020 19935 72076
rect 19935 72020 19964 72076
rect 19980 72020 19991 72076
rect 19991 72020 20044 72076
rect 19900 72016 19964 72020
rect 19980 72016 20044 72020
rect 20060 72016 20124 72080
rect 20140 72016 20204 72080
rect 20220 72016 20284 72080
rect 25740 72076 25804 72080
rect 25740 72020 25771 72076
rect 25771 72020 25804 72076
rect 25740 72016 25804 72020
rect 25820 72016 25884 72080
rect 25900 72016 25964 72080
rect 25980 72016 26044 72080
rect 26060 72016 26124 72080
rect 26140 72016 26204 72080
rect 26220 72016 26284 72080
rect 31740 72016 31804 72080
rect 31820 72016 31884 72080
rect 31900 72016 31964 72080
rect 31980 72016 32044 72080
rect 32060 72016 32124 72080
rect 32140 72016 32204 72080
rect 32220 72016 32284 72080
rect 37740 72016 37804 72080
rect 37820 72016 37884 72080
rect 37900 72016 37964 72080
rect 37980 72016 38044 72080
rect 38060 72016 38124 72080
rect 38140 72016 38204 72080
rect 38220 72016 38284 72080
rect 43740 72016 43804 72080
rect 43820 72016 43884 72080
rect 43900 72016 43964 72080
rect 43980 72016 44044 72080
rect 44060 72016 44124 72080
rect 44140 72016 44204 72080
rect 44220 72016 44284 72080
rect 49740 72076 49804 72080
rect 49820 72076 49884 72080
rect 49740 72020 49754 72076
rect 49754 72020 49804 72076
rect 49820 72020 49834 72076
rect 49834 72020 49884 72076
rect 49740 72016 49804 72020
rect 49820 72016 49884 72020
rect 49900 72016 49964 72080
rect 49980 72016 50044 72080
rect 50060 72016 50124 72080
rect 50140 72016 50204 72080
rect 50220 72016 50284 72080
rect 55740 72016 55804 72080
rect 55820 72016 55884 72080
rect 55900 72016 55964 72080
rect 55980 72016 56044 72080
rect 56060 72016 56124 72080
rect 56140 72016 56204 72080
rect 56220 72016 56284 72080
rect 61740 72016 61804 72080
rect 61820 72016 61884 72080
rect 61900 72016 61964 72080
rect 61980 72016 62044 72080
rect 62060 72016 62124 72080
rect 62140 72016 62204 72080
rect 62220 72016 62284 72080
rect 67740 72016 67804 72080
rect 67820 72016 67884 72080
rect 67900 72016 67964 72080
rect 67980 72016 68044 72080
rect 68060 72016 68124 72080
rect 68140 72016 68204 72080
rect 68220 72016 68284 72080
rect 73740 72016 73804 72080
rect 73820 72016 73884 72080
rect 73900 72016 73964 72080
rect 73980 72016 74044 72080
rect 74060 72016 74124 72080
rect 74140 72016 74204 72080
rect 74220 72016 74284 72080
rect 1740 71936 1804 72000
rect 1820 71936 1884 72000
rect 1900 71936 1964 72000
rect 1980 71936 2044 72000
rect 2060 71936 2124 72000
rect 2140 71936 2204 72000
rect 2220 71996 2284 72000
rect 2220 71940 2276 71996
rect 2276 71940 2284 71996
rect 2220 71936 2284 71940
rect 7740 71936 7804 72000
rect 7820 71936 7884 72000
rect 7900 71936 7964 72000
rect 7980 71936 8044 72000
rect 8060 71936 8124 72000
rect 8140 71936 8204 72000
rect 8220 71936 8284 72000
rect 13740 71936 13804 72000
rect 13820 71936 13884 72000
rect 13900 71936 13964 72000
rect 13980 71936 14044 72000
rect 14060 71936 14124 72000
rect 14140 71996 14204 72000
rect 14140 71940 14155 71996
rect 14155 71940 14204 71996
rect 14140 71936 14204 71940
rect 14220 71936 14284 72000
rect 19740 71936 19804 72000
rect 19820 71936 19884 72000
rect 19900 71996 19964 72000
rect 19980 71996 20044 72000
rect 19900 71940 19935 71996
rect 19935 71940 19964 71996
rect 19980 71940 19991 71996
rect 19991 71940 20044 71996
rect 19900 71936 19964 71940
rect 19980 71936 20044 71940
rect 20060 71936 20124 72000
rect 20140 71936 20204 72000
rect 20220 71936 20284 72000
rect 25740 71996 25804 72000
rect 25740 71940 25771 71996
rect 25771 71940 25804 71996
rect 25740 71936 25804 71940
rect 25820 71936 25884 72000
rect 25900 71936 25964 72000
rect 25980 71936 26044 72000
rect 26060 71936 26124 72000
rect 26140 71936 26204 72000
rect 26220 71936 26284 72000
rect 31740 71936 31804 72000
rect 31820 71936 31884 72000
rect 31900 71936 31964 72000
rect 31980 71936 32044 72000
rect 32060 71936 32124 72000
rect 32140 71936 32204 72000
rect 32220 71936 32284 72000
rect 37740 71936 37804 72000
rect 37820 71936 37884 72000
rect 37900 71936 37964 72000
rect 37980 71936 38044 72000
rect 38060 71936 38124 72000
rect 38140 71936 38204 72000
rect 38220 71936 38284 72000
rect 43740 71936 43804 72000
rect 43820 71936 43884 72000
rect 43900 71936 43964 72000
rect 43980 71936 44044 72000
rect 44060 71936 44124 72000
rect 44140 71936 44204 72000
rect 44220 71936 44284 72000
rect 49740 71996 49804 72000
rect 49820 71996 49884 72000
rect 49740 71940 49754 71996
rect 49754 71940 49804 71996
rect 49820 71940 49834 71996
rect 49834 71940 49884 71996
rect 49740 71936 49804 71940
rect 49820 71936 49884 71940
rect 49900 71936 49964 72000
rect 49980 71936 50044 72000
rect 50060 71936 50124 72000
rect 50140 71936 50204 72000
rect 50220 71936 50284 72000
rect 55740 71936 55804 72000
rect 55820 71936 55884 72000
rect 55900 71936 55964 72000
rect 55980 71936 56044 72000
rect 56060 71936 56124 72000
rect 56140 71936 56204 72000
rect 56220 71936 56284 72000
rect 61740 71936 61804 72000
rect 61820 71936 61884 72000
rect 61900 71936 61964 72000
rect 61980 71936 62044 72000
rect 62060 71936 62124 72000
rect 62140 71936 62204 72000
rect 62220 71936 62284 72000
rect 67740 71936 67804 72000
rect 67820 71936 67884 72000
rect 67900 71936 67964 72000
rect 67980 71936 68044 72000
rect 68060 71936 68124 72000
rect 68140 71936 68204 72000
rect 68220 71936 68284 72000
rect 73740 71936 73804 72000
rect 73820 71936 73884 72000
rect 73900 71936 73964 72000
rect 73980 71936 74044 72000
rect 74060 71936 74124 72000
rect 74140 71936 74204 72000
rect 74220 71936 74284 72000
rect 63540 65240 63604 65244
rect 63540 65184 63554 65240
rect 63554 65184 63604 65240
rect 63540 65180 63604 65184
rect 4740 64528 4804 64592
rect 4820 64528 4884 64592
rect 4900 64528 4964 64592
rect 4980 64528 5044 64592
rect 5060 64528 5124 64592
rect 5140 64528 5204 64592
rect 5220 64528 5284 64592
rect 10740 64528 10804 64592
rect 10820 64528 10884 64592
rect 10900 64528 10964 64592
rect 10980 64528 11044 64592
rect 11060 64528 11124 64592
rect 11140 64528 11204 64592
rect 11220 64528 11284 64592
rect 16740 64528 16804 64592
rect 16820 64528 16884 64592
rect 16900 64528 16964 64592
rect 16980 64528 17044 64592
rect 17060 64528 17124 64592
rect 17140 64588 17204 64592
rect 17220 64588 17284 64592
rect 17140 64532 17192 64588
rect 17192 64532 17204 64588
rect 17220 64532 17248 64588
rect 17248 64532 17284 64588
rect 17140 64528 17204 64532
rect 17220 64528 17284 64532
rect 22740 64528 22804 64592
rect 22820 64528 22884 64592
rect 22900 64528 22964 64592
rect 22980 64588 23044 64592
rect 22980 64532 23028 64588
rect 23028 64532 23044 64588
rect 22980 64528 23044 64532
rect 23060 64528 23124 64592
rect 23140 64528 23204 64592
rect 23220 64528 23284 64592
rect 28740 64588 28804 64592
rect 28740 64532 28752 64588
rect 28752 64532 28804 64588
rect 28740 64528 28804 64532
rect 28820 64528 28884 64592
rect 28900 64528 28964 64592
rect 28980 64528 29044 64592
rect 29060 64528 29124 64592
rect 29140 64528 29204 64592
rect 29220 64528 29284 64592
rect 34740 64528 34804 64592
rect 34820 64528 34884 64592
rect 34900 64528 34964 64592
rect 34980 64528 35044 64592
rect 35060 64528 35124 64592
rect 35140 64528 35204 64592
rect 35220 64528 35284 64592
rect 40740 64528 40804 64592
rect 40820 64528 40884 64592
rect 40900 64528 40964 64592
rect 40980 64528 41044 64592
rect 41060 64528 41124 64592
rect 41140 64528 41204 64592
rect 41220 64528 41284 64592
rect 46740 64528 46804 64592
rect 46820 64528 46884 64592
rect 46900 64528 46964 64592
rect 46980 64528 47044 64592
rect 47060 64528 47124 64592
rect 47140 64528 47204 64592
rect 47220 64528 47284 64592
rect 52740 64528 52804 64592
rect 52820 64528 52884 64592
rect 52900 64528 52964 64592
rect 52980 64528 53044 64592
rect 53060 64528 53124 64592
rect 53140 64528 53204 64592
rect 53220 64528 53284 64592
rect 58740 64528 58804 64592
rect 58820 64528 58884 64592
rect 58900 64528 58964 64592
rect 58980 64528 59044 64592
rect 59060 64528 59124 64592
rect 59140 64588 59204 64592
rect 59140 64532 59196 64588
rect 59196 64532 59204 64588
rect 59140 64528 59204 64532
rect 59220 64528 59284 64592
rect 64740 64528 64804 64592
rect 64820 64528 64884 64592
rect 64900 64528 64964 64592
rect 64980 64528 65044 64592
rect 65060 64528 65124 64592
rect 65140 64528 65204 64592
rect 65220 64528 65284 64592
rect 70740 64528 70804 64592
rect 70820 64528 70884 64592
rect 70900 64528 70964 64592
rect 70980 64528 71044 64592
rect 71060 64528 71124 64592
rect 71140 64528 71204 64592
rect 71220 64528 71284 64592
rect 4740 64448 4804 64512
rect 4820 64448 4884 64512
rect 4900 64448 4964 64512
rect 4980 64448 5044 64512
rect 5060 64448 5124 64512
rect 5140 64448 5204 64512
rect 5220 64448 5284 64512
rect 10740 64448 10804 64512
rect 10820 64448 10884 64512
rect 10900 64448 10964 64512
rect 10980 64448 11044 64512
rect 11060 64448 11124 64512
rect 11140 64448 11204 64512
rect 11220 64448 11284 64512
rect 16740 64448 16804 64512
rect 16820 64448 16884 64512
rect 16900 64448 16964 64512
rect 16980 64448 17044 64512
rect 17060 64448 17124 64512
rect 17140 64508 17204 64512
rect 17220 64508 17284 64512
rect 17140 64452 17192 64508
rect 17192 64452 17204 64508
rect 17220 64452 17248 64508
rect 17248 64452 17284 64508
rect 17140 64448 17204 64452
rect 17220 64448 17284 64452
rect 22740 64448 22804 64512
rect 22820 64448 22884 64512
rect 22900 64448 22964 64512
rect 22980 64508 23044 64512
rect 22980 64452 23028 64508
rect 23028 64452 23044 64508
rect 22980 64448 23044 64452
rect 23060 64448 23124 64512
rect 23140 64448 23204 64512
rect 23220 64448 23284 64512
rect 28740 64508 28804 64512
rect 28740 64452 28752 64508
rect 28752 64452 28804 64508
rect 28740 64448 28804 64452
rect 28820 64448 28884 64512
rect 28900 64448 28964 64512
rect 28980 64448 29044 64512
rect 29060 64448 29124 64512
rect 29140 64448 29204 64512
rect 29220 64448 29284 64512
rect 34740 64448 34804 64512
rect 34820 64448 34884 64512
rect 34900 64448 34964 64512
rect 34980 64448 35044 64512
rect 35060 64448 35124 64512
rect 35140 64448 35204 64512
rect 35220 64448 35284 64512
rect 40740 64448 40804 64512
rect 40820 64448 40884 64512
rect 40900 64448 40964 64512
rect 40980 64448 41044 64512
rect 41060 64448 41124 64512
rect 41140 64448 41204 64512
rect 41220 64448 41284 64512
rect 46740 64448 46804 64512
rect 46820 64448 46884 64512
rect 46900 64448 46964 64512
rect 46980 64448 47044 64512
rect 47060 64448 47124 64512
rect 47140 64448 47204 64512
rect 47220 64448 47284 64512
rect 52740 64448 52804 64512
rect 52820 64448 52884 64512
rect 52900 64448 52964 64512
rect 52980 64448 53044 64512
rect 53060 64448 53124 64512
rect 53140 64448 53204 64512
rect 53220 64448 53284 64512
rect 58740 64448 58804 64512
rect 58820 64448 58884 64512
rect 58900 64448 58964 64512
rect 58980 64448 59044 64512
rect 59060 64448 59124 64512
rect 59140 64508 59204 64512
rect 59140 64452 59196 64508
rect 59196 64452 59204 64508
rect 59140 64448 59204 64452
rect 59220 64448 59284 64512
rect 64740 64448 64804 64512
rect 64820 64448 64884 64512
rect 64900 64448 64964 64512
rect 64980 64448 65044 64512
rect 65060 64448 65124 64512
rect 65140 64448 65204 64512
rect 65220 64448 65284 64512
rect 70740 64448 70804 64512
rect 70820 64448 70884 64512
rect 70900 64448 70964 64512
rect 70980 64448 71044 64512
rect 71060 64448 71124 64512
rect 71140 64448 71204 64512
rect 71220 64448 71284 64512
rect 4740 64368 4804 64432
rect 4820 64368 4884 64432
rect 4900 64368 4964 64432
rect 4980 64368 5044 64432
rect 5060 64368 5124 64432
rect 5140 64368 5204 64432
rect 5220 64368 5284 64432
rect 10740 64368 10804 64432
rect 10820 64368 10884 64432
rect 10900 64368 10964 64432
rect 10980 64368 11044 64432
rect 11060 64368 11124 64432
rect 11140 64368 11204 64432
rect 11220 64368 11284 64432
rect 16740 64368 16804 64432
rect 16820 64368 16884 64432
rect 16900 64368 16964 64432
rect 16980 64368 17044 64432
rect 17060 64368 17124 64432
rect 17140 64428 17204 64432
rect 17220 64428 17284 64432
rect 17140 64372 17192 64428
rect 17192 64372 17204 64428
rect 17220 64372 17248 64428
rect 17248 64372 17284 64428
rect 17140 64368 17204 64372
rect 17220 64368 17284 64372
rect 22740 64368 22804 64432
rect 22820 64368 22884 64432
rect 22900 64368 22964 64432
rect 22980 64428 23044 64432
rect 22980 64372 23028 64428
rect 23028 64372 23044 64428
rect 22980 64368 23044 64372
rect 23060 64368 23124 64432
rect 23140 64368 23204 64432
rect 23220 64368 23284 64432
rect 28740 64428 28804 64432
rect 28740 64372 28752 64428
rect 28752 64372 28804 64428
rect 28740 64368 28804 64372
rect 28820 64368 28884 64432
rect 28900 64368 28964 64432
rect 28980 64368 29044 64432
rect 29060 64368 29124 64432
rect 29140 64368 29204 64432
rect 29220 64368 29284 64432
rect 34740 64368 34804 64432
rect 34820 64368 34884 64432
rect 34900 64368 34964 64432
rect 34980 64368 35044 64432
rect 35060 64368 35124 64432
rect 35140 64368 35204 64432
rect 35220 64368 35284 64432
rect 40740 64368 40804 64432
rect 40820 64368 40884 64432
rect 40900 64368 40964 64432
rect 40980 64368 41044 64432
rect 41060 64368 41124 64432
rect 41140 64368 41204 64432
rect 41220 64368 41284 64432
rect 46740 64368 46804 64432
rect 46820 64368 46884 64432
rect 46900 64368 46964 64432
rect 46980 64368 47044 64432
rect 47060 64368 47124 64432
rect 47140 64368 47204 64432
rect 47220 64368 47284 64432
rect 52740 64368 52804 64432
rect 52820 64368 52884 64432
rect 52900 64368 52964 64432
rect 52980 64368 53044 64432
rect 53060 64368 53124 64432
rect 53140 64368 53204 64432
rect 53220 64368 53284 64432
rect 58740 64368 58804 64432
rect 58820 64368 58884 64432
rect 58900 64368 58964 64432
rect 58980 64368 59044 64432
rect 59060 64368 59124 64432
rect 59140 64428 59204 64432
rect 59140 64372 59196 64428
rect 59196 64372 59204 64428
rect 59140 64368 59204 64372
rect 59220 64368 59284 64432
rect 64740 64368 64804 64432
rect 64820 64368 64884 64432
rect 64900 64368 64964 64432
rect 64980 64368 65044 64432
rect 65060 64368 65124 64432
rect 65140 64368 65204 64432
rect 65220 64368 65284 64432
rect 70740 64368 70804 64432
rect 70820 64368 70884 64432
rect 70900 64368 70964 64432
rect 70980 64368 71044 64432
rect 71060 64368 71124 64432
rect 71140 64368 71204 64432
rect 71220 64368 71284 64432
rect 4740 64288 4804 64352
rect 4820 64288 4884 64352
rect 4900 64288 4964 64352
rect 4980 64288 5044 64352
rect 5060 64288 5124 64352
rect 5140 64288 5204 64352
rect 5220 64288 5284 64352
rect 10740 64288 10804 64352
rect 10820 64288 10884 64352
rect 10900 64288 10964 64352
rect 10980 64288 11044 64352
rect 11060 64288 11124 64352
rect 11140 64288 11204 64352
rect 11220 64288 11284 64352
rect 16740 64288 16804 64352
rect 16820 64288 16884 64352
rect 16900 64288 16964 64352
rect 16980 64288 17044 64352
rect 17060 64288 17124 64352
rect 17140 64348 17204 64352
rect 17220 64348 17284 64352
rect 17140 64292 17192 64348
rect 17192 64292 17204 64348
rect 17220 64292 17248 64348
rect 17248 64292 17284 64348
rect 17140 64288 17204 64292
rect 17220 64288 17284 64292
rect 22740 64288 22804 64352
rect 22820 64288 22884 64352
rect 22900 64288 22964 64352
rect 22980 64348 23044 64352
rect 22980 64292 23028 64348
rect 23028 64292 23044 64348
rect 22980 64288 23044 64292
rect 23060 64288 23124 64352
rect 23140 64288 23204 64352
rect 23220 64288 23284 64352
rect 28740 64348 28804 64352
rect 28740 64292 28752 64348
rect 28752 64292 28804 64348
rect 28740 64288 28804 64292
rect 28820 64288 28884 64352
rect 28900 64288 28964 64352
rect 28980 64288 29044 64352
rect 29060 64288 29124 64352
rect 29140 64288 29204 64352
rect 29220 64288 29284 64352
rect 34740 64288 34804 64352
rect 34820 64288 34884 64352
rect 34900 64288 34964 64352
rect 34980 64288 35044 64352
rect 35060 64288 35124 64352
rect 35140 64288 35204 64352
rect 35220 64288 35284 64352
rect 40740 64288 40804 64352
rect 40820 64288 40884 64352
rect 40900 64288 40964 64352
rect 40980 64288 41044 64352
rect 41060 64288 41124 64352
rect 41140 64288 41204 64352
rect 41220 64288 41284 64352
rect 46740 64288 46804 64352
rect 46820 64288 46884 64352
rect 46900 64288 46964 64352
rect 46980 64288 47044 64352
rect 47060 64288 47124 64352
rect 47140 64288 47204 64352
rect 47220 64288 47284 64352
rect 52740 64288 52804 64352
rect 52820 64288 52884 64352
rect 52900 64288 52964 64352
rect 52980 64288 53044 64352
rect 53060 64288 53124 64352
rect 53140 64288 53204 64352
rect 53220 64288 53284 64352
rect 58740 64288 58804 64352
rect 58820 64288 58884 64352
rect 58900 64288 58964 64352
rect 58980 64288 59044 64352
rect 59060 64288 59124 64352
rect 59140 64348 59204 64352
rect 59140 64292 59196 64348
rect 59196 64292 59204 64348
rect 59140 64288 59204 64292
rect 59220 64288 59284 64352
rect 64740 64288 64804 64352
rect 64820 64288 64884 64352
rect 64900 64288 64964 64352
rect 64980 64288 65044 64352
rect 65060 64288 65124 64352
rect 65140 64288 65204 64352
rect 65220 64288 65284 64352
rect 70740 64288 70804 64352
rect 70820 64288 70884 64352
rect 70900 64288 70964 64352
rect 70980 64288 71044 64352
rect 71060 64288 71124 64352
rect 71140 64288 71204 64352
rect 71220 64288 71284 64352
rect 63724 63140 63788 63204
rect 1740 62176 1804 62240
rect 1820 62176 1884 62240
rect 1900 62176 1964 62240
rect 1980 62176 2044 62240
rect 2060 62176 2124 62240
rect 2140 62176 2204 62240
rect 2220 62236 2284 62240
rect 2220 62180 2276 62236
rect 2276 62180 2284 62236
rect 2220 62176 2284 62180
rect 7740 62176 7804 62240
rect 7820 62176 7884 62240
rect 7900 62176 7964 62240
rect 7980 62176 8044 62240
rect 8060 62176 8124 62240
rect 8140 62176 8204 62240
rect 8220 62176 8284 62240
rect 13740 62176 13804 62240
rect 13820 62176 13884 62240
rect 13900 62176 13964 62240
rect 13980 62176 14044 62240
rect 14060 62176 14124 62240
rect 14140 62236 14204 62240
rect 14140 62180 14155 62236
rect 14155 62180 14204 62236
rect 14140 62176 14204 62180
rect 14220 62176 14284 62240
rect 19740 62176 19804 62240
rect 19820 62176 19884 62240
rect 19900 62236 19964 62240
rect 19980 62236 20044 62240
rect 19900 62180 19935 62236
rect 19935 62180 19964 62236
rect 19980 62180 19991 62236
rect 19991 62180 20044 62236
rect 19900 62176 19964 62180
rect 19980 62176 20044 62180
rect 20060 62176 20124 62240
rect 20140 62176 20204 62240
rect 20220 62176 20284 62240
rect 25740 62236 25804 62240
rect 25740 62180 25771 62236
rect 25771 62180 25804 62236
rect 25740 62176 25804 62180
rect 25820 62176 25884 62240
rect 25900 62176 25964 62240
rect 25980 62176 26044 62240
rect 26060 62176 26124 62240
rect 26140 62176 26204 62240
rect 26220 62176 26284 62240
rect 31740 62176 31804 62240
rect 31820 62176 31884 62240
rect 31900 62176 31964 62240
rect 31980 62176 32044 62240
rect 32060 62176 32124 62240
rect 32140 62176 32204 62240
rect 32220 62176 32284 62240
rect 37740 62176 37804 62240
rect 37820 62176 37884 62240
rect 37900 62176 37964 62240
rect 37980 62176 38044 62240
rect 38060 62176 38124 62240
rect 38140 62176 38204 62240
rect 38220 62176 38284 62240
rect 43740 62176 43804 62240
rect 43820 62176 43884 62240
rect 43900 62176 43964 62240
rect 43980 62176 44044 62240
rect 44060 62176 44124 62240
rect 44140 62176 44204 62240
rect 44220 62176 44284 62240
rect 49740 62236 49804 62240
rect 49820 62236 49884 62240
rect 49740 62180 49754 62236
rect 49754 62180 49804 62236
rect 49820 62180 49834 62236
rect 49834 62180 49884 62236
rect 49740 62176 49804 62180
rect 49820 62176 49884 62180
rect 49900 62176 49964 62240
rect 49980 62176 50044 62240
rect 50060 62176 50124 62240
rect 50140 62176 50204 62240
rect 50220 62176 50284 62240
rect 55740 62176 55804 62240
rect 55820 62176 55884 62240
rect 55900 62176 55964 62240
rect 55980 62176 56044 62240
rect 56060 62176 56124 62240
rect 56140 62176 56204 62240
rect 56220 62176 56284 62240
rect 61740 62176 61804 62240
rect 61820 62176 61884 62240
rect 61900 62176 61964 62240
rect 61980 62176 62044 62240
rect 62060 62176 62124 62240
rect 62140 62176 62204 62240
rect 62220 62176 62284 62240
rect 67740 62176 67804 62240
rect 67820 62176 67884 62240
rect 67900 62176 67964 62240
rect 67980 62176 68044 62240
rect 68060 62176 68124 62240
rect 68140 62176 68204 62240
rect 68220 62176 68284 62240
rect 73740 62176 73804 62240
rect 73820 62176 73884 62240
rect 73900 62176 73964 62240
rect 73980 62176 74044 62240
rect 74060 62176 74124 62240
rect 74140 62176 74204 62240
rect 74220 62176 74284 62240
rect 1740 62096 1804 62160
rect 1820 62096 1884 62160
rect 1900 62096 1964 62160
rect 1980 62096 2044 62160
rect 2060 62096 2124 62160
rect 2140 62096 2204 62160
rect 2220 62156 2284 62160
rect 2220 62100 2276 62156
rect 2276 62100 2284 62156
rect 2220 62096 2284 62100
rect 7740 62096 7804 62160
rect 7820 62096 7884 62160
rect 7900 62096 7964 62160
rect 7980 62096 8044 62160
rect 8060 62096 8124 62160
rect 8140 62096 8204 62160
rect 8220 62096 8284 62160
rect 13740 62096 13804 62160
rect 13820 62096 13884 62160
rect 13900 62096 13964 62160
rect 13980 62096 14044 62160
rect 14060 62096 14124 62160
rect 14140 62156 14204 62160
rect 14140 62100 14155 62156
rect 14155 62100 14204 62156
rect 14140 62096 14204 62100
rect 14220 62096 14284 62160
rect 19740 62096 19804 62160
rect 19820 62096 19884 62160
rect 19900 62156 19964 62160
rect 19980 62156 20044 62160
rect 19900 62100 19935 62156
rect 19935 62100 19964 62156
rect 19980 62100 19991 62156
rect 19991 62100 20044 62156
rect 19900 62096 19964 62100
rect 19980 62096 20044 62100
rect 20060 62096 20124 62160
rect 20140 62096 20204 62160
rect 20220 62096 20284 62160
rect 25740 62156 25804 62160
rect 25740 62100 25771 62156
rect 25771 62100 25804 62156
rect 25740 62096 25804 62100
rect 25820 62096 25884 62160
rect 25900 62096 25964 62160
rect 25980 62096 26044 62160
rect 26060 62096 26124 62160
rect 26140 62096 26204 62160
rect 26220 62096 26284 62160
rect 31740 62096 31804 62160
rect 31820 62096 31884 62160
rect 31900 62096 31964 62160
rect 31980 62096 32044 62160
rect 32060 62096 32124 62160
rect 32140 62096 32204 62160
rect 32220 62096 32284 62160
rect 37740 62096 37804 62160
rect 37820 62096 37884 62160
rect 37900 62096 37964 62160
rect 37980 62096 38044 62160
rect 38060 62096 38124 62160
rect 38140 62096 38204 62160
rect 38220 62096 38284 62160
rect 43740 62096 43804 62160
rect 43820 62096 43884 62160
rect 43900 62096 43964 62160
rect 43980 62096 44044 62160
rect 44060 62096 44124 62160
rect 44140 62096 44204 62160
rect 44220 62096 44284 62160
rect 49740 62156 49804 62160
rect 49820 62156 49884 62160
rect 49740 62100 49754 62156
rect 49754 62100 49804 62156
rect 49820 62100 49834 62156
rect 49834 62100 49884 62156
rect 49740 62096 49804 62100
rect 49820 62096 49884 62100
rect 49900 62096 49964 62160
rect 49980 62096 50044 62160
rect 50060 62096 50124 62160
rect 50140 62096 50204 62160
rect 50220 62096 50284 62160
rect 55740 62096 55804 62160
rect 55820 62096 55884 62160
rect 55900 62096 55964 62160
rect 55980 62096 56044 62160
rect 56060 62096 56124 62160
rect 56140 62096 56204 62160
rect 56220 62096 56284 62160
rect 61740 62096 61804 62160
rect 61820 62096 61884 62160
rect 61900 62096 61964 62160
rect 61980 62096 62044 62160
rect 62060 62096 62124 62160
rect 62140 62096 62204 62160
rect 62220 62096 62284 62160
rect 67740 62096 67804 62160
rect 67820 62096 67884 62160
rect 67900 62096 67964 62160
rect 67980 62096 68044 62160
rect 68060 62096 68124 62160
rect 68140 62096 68204 62160
rect 68220 62096 68284 62160
rect 73740 62096 73804 62160
rect 73820 62096 73884 62160
rect 73900 62096 73964 62160
rect 73980 62096 74044 62160
rect 74060 62096 74124 62160
rect 74140 62096 74204 62160
rect 74220 62096 74284 62160
rect 1740 62016 1804 62080
rect 1820 62016 1884 62080
rect 1900 62016 1964 62080
rect 1980 62016 2044 62080
rect 2060 62016 2124 62080
rect 2140 62016 2204 62080
rect 2220 62076 2284 62080
rect 2220 62020 2276 62076
rect 2276 62020 2284 62076
rect 2220 62016 2284 62020
rect 7740 62016 7804 62080
rect 7820 62016 7884 62080
rect 7900 62016 7964 62080
rect 7980 62016 8044 62080
rect 8060 62016 8124 62080
rect 8140 62016 8204 62080
rect 8220 62016 8284 62080
rect 13740 62016 13804 62080
rect 13820 62016 13884 62080
rect 13900 62016 13964 62080
rect 13980 62016 14044 62080
rect 14060 62016 14124 62080
rect 14140 62076 14204 62080
rect 14140 62020 14155 62076
rect 14155 62020 14204 62076
rect 14140 62016 14204 62020
rect 14220 62016 14284 62080
rect 19740 62016 19804 62080
rect 19820 62016 19884 62080
rect 19900 62076 19964 62080
rect 19980 62076 20044 62080
rect 19900 62020 19935 62076
rect 19935 62020 19964 62076
rect 19980 62020 19991 62076
rect 19991 62020 20044 62076
rect 19900 62016 19964 62020
rect 19980 62016 20044 62020
rect 20060 62016 20124 62080
rect 20140 62016 20204 62080
rect 20220 62016 20284 62080
rect 25740 62076 25804 62080
rect 25740 62020 25771 62076
rect 25771 62020 25804 62076
rect 25740 62016 25804 62020
rect 25820 62016 25884 62080
rect 25900 62016 25964 62080
rect 25980 62016 26044 62080
rect 26060 62016 26124 62080
rect 26140 62016 26204 62080
rect 26220 62016 26284 62080
rect 31740 62016 31804 62080
rect 31820 62016 31884 62080
rect 31900 62016 31964 62080
rect 31980 62016 32044 62080
rect 32060 62016 32124 62080
rect 32140 62016 32204 62080
rect 32220 62016 32284 62080
rect 37740 62016 37804 62080
rect 37820 62016 37884 62080
rect 37900 62016 37964 62080
rect 37980 62016 38044 62080
rect 38060 62016 38124 62080
rect 38140 62016 38204 62080
rect 38220 62016 38284 62080
rect 43740 62016 43804 62080
rect 43820 62016 43884 62080
rect 43900 62016 43964 62080
rect 43980 62016 44044 62080
rect 44060 62016 44124 62080
rect 44140 62016 44204 62080
rect 44220 62016 44284 62080
rect 49740 62076 49804 62080
rect 49820 62076 49884 62080
rect 49740 62020 49754 62076
rect 49754 62020 49804 62076
rect 49820 62020 49834 62076
rect 49834 62020 49884 62076
rect 49740 62016 49804 62020
rect 49820 62016 49884 62020
rect 49900 62016 49964 62080
rect 49980 62016 50044 62080
rect 50060 62016 50124 62080
rect 50140 62016 50204 62080
rect 50220 62016 50284 62080
rect 55740 62016 55804 62080
rect 55820 62016 55884 62080
rect 55900 62016 55964 62080
rect 55980 62016 56044 62080
rect 56060 62016 56124 62080
rect 56140 62016 56204 62080
rect 56220 62016 56284 62080
rect 61740 62016 61804 62080
rect 61820 62016 61884 62080
rect 61900 62016 61964 62080
rect 61980 62016 62044 62080
rect 62060 62016 62124 62080
rect 62140 62016 62204 62080
rect 62220 62016 62284 62080
rect 67740 62016 67804 62080
rect 67820 62016 67884 62080
rect 67900 62016 67964 62080
rect 67980 62016 68044 62080
rect 68060 62016 68124 62080
rect 68140 62016 68204 62080
rect 68220 62016 68284 62080
rect 73740 62016 73804 62080
rect 73820 62016 73884 62080
rect 73900 62016 73964 62080
rect 73980 62016 74044 62080
rect 74060 62016 74124 62080
rect 74140 62016 74204 62080
rect 74220 62016 74284 62080
rect 1740 61936 1804 62000
rect 1820 61936 1884 62000
rect 1900 61936 1964 62000
rect 1980 61936 2044 62000
rect 2060 61936 2124 62000
rect 2140 61936 2204 62000
rect 2220 61996 2284 62000
rect 2220 61940 2276 61996
rect 2276 61940 2284 61996
rect 2220 61936 2284 61940
rect 7740 61936 7804 62000
rect 7820 61936 7884 62000
rect 7900 61936 7964 62000
rect 7980 61936 8044 62000
rect 8060 61936 8124 62000
rect 8140 61936 8204 62000
rect 8220 61936 8284 62000
rect 13740 61936 13804 62000
rect 13820 61936 13884 62000
rect 13900 61936 13964 62000
rect 13980 61936 14044 62000
rect 14060 61936 14124 62000
rect 14140 61996 14204 62000
rect 14140 61940 14155 61996
rect 14155 61940 14204 61996
rect 14140 61936 14204 61940
rect 14220 61936 14284 62000
rect 19740 61936 19804 62000
rect 19820 61936 19884 62000
rect 19900 61996 19964 62000
rect 19980 61996 20044 62000
rect 19900 61940 19935 61996
rect 19935 61940 19964 61996
rect 19980 61940 19991 61996
rect 19991 61940 20044 61996
rect 19900 61936 19964 61940
rect 19980 61936 20044 61940
rect 20060 61936 20124 62000
rect 20140 61936 20204 62000
rect 20220 61936 20284 62000
rect 25740 61996 25804 62000
rect 25740 61940 25771 61996
rect 25771 61940 25804 61996
rect 25740 61936 25804 61940
rect 25820 61936 25884 62000
rect 25900 61936 25964 62000
rect 25980 61936 26044 62000
rect 26060 61936 26124 62000
rect 26140 61936 26204 62000
rect 26220 61936 26284 62000
rect 31740 61936 31804 62000
rect 31820 61936 31884 62000
rect 31900 61936 31964 62000
rect 31980 61936 32044 62000
rect 32060 61936 32124 62000
rect 32140 61936 32204 62000
rect 32220 61936 32284 62000
rect 37740 61936 37804 62000
rect 37820 61936 37884 62000
rect 37900 61936 37964 62000
rect 37980 61936 38044 62000
rect 38060 61936 38124 62000
rect 38140 61936 38204 62000
rect 38220 61936 38284 62000
rect 43740 61936 43804 62000
rect 43820 61936 43884 62000
rect 43900 61936 43964 62000
rect 43980 61936 44044 62000
rect 44060 61936 44124 62000
rect 44140 61936 44204 62000
rect 44220 61936 44284 62000
rect 49740 61996 49804 62000
rect 49820 61996 49884 62000
rect 49740 61940 49754 61996
rect 49754 61940 49804 61996
rect 49820 61940 49834 61996
rect 49834 61940 49884 61996
rect 49740 61936 49804 61940
rect 49820 61936 49884 61940
rect 49900 61936 49964 62000
rect 49980 61936 50044 62000
rect 50060 61936 50124 62000
rect 50140 61936 50204 62000
rect 50220 61936 50284 62000
rect 55740 61936 55804 62000
rect 55820 61936 55884 62000
rect 55900 61936 55964 62000
rect 55980 61936 56044 62000
rect 56060 61936 56124 62000
rect 56140 61936 56204 62000
rect 56220 61936 56284 62000
rect 61740 61936 61804 62000
rect 61820 61936 61884 62000
rect 61900 61936 61964 62000
rect 61980 61936 62044 62000
rect 62060 61936 62124 62000
rect 62140 61936 62204 62000
rect 62220 61936 62284 62000
rect 67740 61936 67804 62000
rect 67820 61936 67884 62000
rect 67900 61936 67964 62000
rect 67980 61936 68044 62000
rect 68060 61936 68124 62000
rect 68140 61936 68204 62000
rect 68220 61936 68284 62000
rect 73740 61936 73804 62000
rect 73820 61936 73884 62000
rect 73900 61936 73964 62000
rect 73980 61936 74044 62000
rect 74060 61936 74124 62000
rect 74140 61936 74204 62000
rect 74220 61936 74284 62000
rect 63908 60964 63972 61028
rect 64092 58652 64156 58716
rect 64276 56612 64340 56676
rect 69060 54708 69124 54772
rect 4740 54528 4804 54592
rect 4820 54528 4884 54592
rect 4900 54528 4964 54592
rect 4980 54528 5044 54592
rect 5060 54528 5124 54592
rect 5140 54528 5204 54592
rect 5220 54528 5284 54592
rect 10740 54528 10804 54592
rect 10820 54528 10884 54592
rect 10900 54528 10964 54592
rect 10980 54528 11044 54592
rect 11060 54528 11124 54592
rect 11140 54528 11204 54592
rect 11220 54528 11284 54592
rect 16740 54528 16804 54592
rect 16820 54528 16884 54592
rect 16900 54528 16964 54592
rect 16980 54528 17044 54592
rect 17060 54528 17124 54592
rect 17140 54588 17204 54592
rect 17220 54588 17284 54592
rect 17140 54532 17192 54588
rect 17192 54532 17204 54588
rect 17220 54532 17248 54588
rect 17248 54532 17284 54588
rect 17140 54528 17204 54532
rect 17220 54528 17284 54532
rect 22740 54528 22804 54592
rect 22820 54528 22884 54592
rect 22900 54528 22964 54592
rect 22980 54588 23044 54592
rect 22980 54532 23028 54588
rect 23028 54532 23044 54588
rect 22980 54528 23044 54532
rect 23060 54528 23124 54592
rect 23140 54528 23204 54592
rect 23220 54528 23284 54592
rect 28740 54588 28804 54592
rect 28740 54532 28752 54588
rect 28752 54532 28804 54588
rect 28740 54528 28804 54532
rect 28820 54528 28884 54592
rect 28900 54528 28964 54592
rect 28980 54528 29044 54592
rect 29060 54528 29124 54592
rect 29140 54528 29204 54592
rect 29220 54528 29284 54592
rect 34740 54528 34804 54592
rect 34820 54528 34884 54592
rect 34900 54528 34964 54592
rect 34980 54528 35044 54592
rect 35060 54528 35124 54592
rect 35140 54528 35204 54592
rect 35220 54528 35284 54592
rect 40740 54528 40804 54592
rect 40820 54528 40884 54592
rect 40900 54528 40964 54592
rect 40980 54528 41044 54592
rect 41060 54528 41124 54592
rect 41140 54528 41204 54592
rect 41220 54528 41284 54592
rect 46740 54528 46804 54592
rect 46820 54528 46884 54592
rect 46900 54528 46964 54592
rect 46980 54528 47044 54592
rect 47060 54528 47124 54592
rect 47140 54528 47204 54592
rect 47220 54528 47284 54592
rect 52740 54528 52804 54592
rect 52820 54528 52884 54592
rect 52900 54528 52964 54592
rect 52980 54528 53044 54592
rect 53060 54528 53124 54592
rect 53140 54528 53204 54592
rect 53220 54528 53284 54592
rect 58740 54528 58804 54592
rect 58820 54528 58884 54592
rect 58900 54528 58964 54592
rect 58980 54528 59044 54592
rect 59060 54528 59124 54592
rect 59140 54588 59204 54592
rect 59140 54532 59196 54588
rect 59196 54532 59204 54588
rect 59140 54528 59204 54532
rect 59220 54528 59284 54592
rect 64740 54528 64804 54592
rect 64820 54528 64884 54592
rect 64900 54528 64964 54592
rect 64980 54528 65044 54592
rect 65060 54528 65124 54592
rect 65140 54528 65204 54592
rect 65220 54528 65284 54592
rect 70740 54528 70804 54592
rect 70820 54528 70884 54592
rect 70900 54528 70964 54592
rect 70980 54528 71044 54592
rect 71060 54528 71124 54592
rect 71140 54528 71204 54592
rect 71220 54528 71284 54592
rect 4740 54448 4804 54512
rect 4820 54448 4884 54512
rect 4900 54448 4964 54512
rect 4980 54448 5044 54512
rect 5060 54448 5124 54512
rect 5140 54448 5204 54512
rect 5220 54448 5284 54512
rect 10740 54448 10804 54512
rect 10820 54448 10884 54512
rect 10900 54448 10964 54512
rect 10980 54448 11044 54512
rect 11060 54448 11124 54512
rect 11140 54448 11204 54512
rect 11220 54448 11284 54512
rect 16740 54448 16804 54512
rect 16820 54448 16884 54512
rect 16900 54448 16964 54512
rect 16980 54448 17044 54512
rect 17060 54448 17124 54512
rect 17140 54508 17204 54512
rect 17220 54508 17284 54512
rect 17140 54452 17192 54508
rect 17192 54452 17204 54508
rect 17220 54452 17248 54508
rect 17248 54452 17284 54508
rect 17140 54448 17204 54452
rect 17220 54448 17284 54452
rect 22740 54448 22804 54512
rect 22820 54448 22884 54512
rect 22900 54448 22964 54512
rect 22980 54508 23044 54512
rect 22980 54452 23028 54508
rect 23028 54452 23044 54508
rect 22980 54448 23044 54452
rect 23060 54448 23124 54512
rect 23140 54448 23204 54512
rect 23220 54448 23284 54512
rect 28740 54508 28804 54512
rect 28740 54452 28752 54508
rect 28752 54452 28804 54508
rect 28740 54448 28804 54452
rect 28820 54448 28884 54512
rect 28900 54448 28964 54512
rect 28980 54448 29044 54512
rect 29060 54448 29124 54512
rect 29140 54448 29204 54512
rect 29220 54448 29284 54512
rect 34740 54448 34804 54512
rect 34820 54448 34884 54512
rect 34900 54448 34964 54512
rect 34980 54448 35044 54512
rect 35060 54448 35124 54512
rect 35140 54448 35204 54512
rect 35220 54448 35284 54512
rect 40740 54448 40804 54512
rect 40820 54448 40884 54512
rect 40900 54448 40964 54512
rect 40980 54448 41044 54512
rect 41060 54448 41124 54512
rect 41140 54448 41204 54512
rect 41220 54448 41284 54512
rect 46740 54448 46804 54512
rect 46820 54448 46884 54512
rect 46900 54448 46964 54512
rect 46980 54448 47044 54512
rect 47060 54448 47124 54512
rect 47140 54448 47204 54512
rect 47220 54448 47284 54512
rect 52740 54448 52804 54512
rect 52820 54448 52884 54512
rect 52900 54448 52964 54512
rect 52980 54448 53044 54512
rect 53060 54448 53124 54512
rect 53140 54448 53204 54512
rect 53220 54448 53284 54512
rect 58740 54448 58804 54512
rect 58820 54448 58884 54512
rect 58900 54448 58964 54512
rect 58980 54448 59044 54512
rect 59060 54448 59124 54512
rect 59140 54508 59204 54512
rect 59140 54452 59196 54508
rect 59196 54452 59204 54508
rect 59140 54448 59204 54452
rect 59220 54448 59284 54512
rect 64740 54448 64804 54512
rect 64820 54448 64884 54512
rect 64900 54448 64964 54512
rect 64980 54448 65044 54512
rect 65060 54448 65124 54512
rect 65140 54448 65204 54512
rect 65220 54448 65284 54512
rect 70740 54448 70804 54512
rect 70820 54448 70884 54512
rect 70900 54448 70964 54512
rect 70980 54448 71044 54512
rect 71060 54448 71124 54512
rect 71140 54448 71204 54512
rect 71220 54448 71284 54512
rect 4740 54368 4804 54432
rect 4820 54368 4884 54432
rect 4900 54368 4964 54432
rect 4980 54368 5044 54432
rect 5060 54368 5124 54432
rect 5140 54368 5204 54432
rect 5220 54368 5284 54432
rect 10740 54368 10804 54432
rect 10820 54368 10884 54432
rect 10900 54368 10964 54432
rect 10980 54368 11044 54432
rect 11060 54368 11124 54432
rect 11140 54368 11204 54432
rect 11220 54368 11284 54432
rect 16740 54368 16804 54432
rect 16820 54368 16884 54432
rect 16900 54368 16964 54432
rect 16980 54368 17044 54432
rect 17060 54368 17124 54432
rect 17140 54428 17204 54432
rect 17220 54428 17284 54432
rect 17140 54372 17192 54428
rect 17192 54372 17204 54428
rect 17220 54372 17248 54428
rect 17248 54372 17284 54428
rect 17140 54368 17204 54372
rect 17220 54368 17284 54372
rect 22740 54368 22804 54432
rect 22820 54368 22884 54432
rect 22900 54368 22964 54432
rect 22980 54428 23044 54432
rect 22980 54372 23028 54428
rect 23028 54372 23044 54428
rect 22980 54368 23044 54372
rect 23060 54368 23124 54432
rect 23140 54368 23204 54432
rect 23220 54368 23284 54432
rect 28740 54428 28804 54432
rect 28740 54372 28752 54428
rect 28752 54372 28804 54428
rect 28740 54368 28804 54372
rect 28820 54368 28884 54432
rect 28900 54368 28964 54432
rect 28980 54368 29044 54432
rect 29060 54368 29124 54432
rect 29140 54368 29204 54432
rect 29220 54368 29284 54432
rect 34740 54368 34804 54432
rect 34820 54368 34884 54432
rect 34900 54368 34964 54432
rect 34980 54368 35044 54432
rect 35060 54368 35124 54432
rect 35140 54368 35204 54432
rect 35220 54368 35284 54432
rect 40740 54368 40804 54432
rect 40820 54368 40884 54432
rect 40900 54368 40964 54432
rect 40980 54368 41044 54432
rect 41060 54368 41124 54432
rect 41140 54368 41204 54432
rect 41220 54368 41284 54432
rect 46740 54368 46804 54432
rect 46820 54368 46884 54432
rect 46900 54368 46964 54432
rect 46980 54368 47044 54432
rect 47060 54368 47124 54432
rect 47140 54368 47204 54432
rect 47220 54368 47284 54432
rect 52740 54368 52804 54432
rect 52820 54368 52884 54432
rect 52900 54368 52964 54432
rect 52980 54368 53044 54432
rect 53060 54368 53124 54432
rect 53140 54368 53204 54432
rect 53220 54368 53284 54432
rect 58740 54368 58804 54432
rect 58820 54368 58884 54432
rect 58900 54368 58964 54432
rect 58980 54368 59044 54432
rect 59060 54368 59124 54432
rect 59140 54428 59204 54432
rect 59140 54372 59196 54428
rect 59196 54372 59204 54428
rect 59140 54368 59204 54372
rect 59220 54368 59284 54432
rect 64740 54368 64804 54432
rect 64820 54368 64884 54432
rect 64900 54368 64964 54432
rect 64980 54368 65044 54432
rect 65060 54368 65124 54432
rect 65140 54368 65204 54432
rect 65220 54368 65284 54432
rect 70740 54368 70804 54432
rect 70820 54368 70884 54432
rect 70900 54368 70964 54432
rect 70980 54368 71044 54432
rect 71060 54368 71124 54432
rect 71140 54368 71204 54432
rect 71220 54368 71284 54432
rect 4740 54288 4804 54352
rect 4820 54288 4884 54352
rect 4900 54288 4964 54352
rect 4980 54288 5044 54352
rect 5060 54288 5124 54352
rect 5140 54288 5204 54352
rect 5220 54288 5284 54352
rect 10740 54288 10804 54352
rect 10820 54288 10884 54352
rect 10900 54288 10964 54352
rect 10980 54288 11044 54352
rect 11060 54288 11124 54352
rect 11140 54288 11204 54352
rect 11220 54288 11284 54352
rect 16740 54288 16804 54352
rect 16820 54288 16884 54352
rect 16900 54288 16964 54352
rect 16980 54288 17044 54352
rect 17060 54288 17124 54352
rect 17140 54348 17204 54352
rect 17220 54348 17284 54352
rect 17140 54292 17192 54348
rect 17192 54292 17204 54348
rect 17220 54292 17248 54348
rect 17248 54292 17284 54348
rect 17140 54288 17204 54292
rect 17220 54288 17284 54292
rect 22740 54288 22804 54352
rect 22820 54288 22884 54352
rect 22900 54288 22964 54352
rect 22980 54348 23044 54352
rect 22980 54292 23028 54348
rect 23028 54292 23044 54348
rect 22980 54288 23044 54292
rect 23060 54288 23124 54352
rect 23140 54288 23204 54352
rect 23220 54288 23284 54352
rect 28740 54348 28804 54352
rect 28740 54292 28752 54348
rect 28752 54292 28804 54348
rect 28740 54288 28804 54292
rect 28820 54288 28884 54352
rect 28900 54288 28964 54352
rect 28980 54288 29044 54352
rect 29060 54288 29124 54352
rect 29140 54288 29204 54352
rect 29220 54288 29284 54352
rect 34740 54288 34804 54352
rect 34820 54288 34884 54352
rect 34900 54288 34964 54352
rect 34980 54288 35044 54352
rect 35060 54288 35124 54352
rect 35140 54288 35204 54352
rect 35220 54288 35284 54352
rect 40740 54288 40804 54352
rect 40820 54288 40884 54352
rect 40900 54288 40964 54352
rect 40980 54288 41044 54352
rect 41060 54288 41124 54352
rect 41140 54288 41204 54352
rect 41220 54288 41284 54352
rect 46740 54288 46804 54352
rect 46820 54288 46884 54352
rect 46900 54288 46964 54352
rect 46980 54288 47044 54352
rect 47060 54288 47124 54352
rect 47140 54288 47204 54352
rect 47220 54288 47284 54352
rect 52740 54288 52804 54352
rect 52820 54288 52884 54352
rect 52900 54288 52964 54352
rect 52980 54288 53044 54352
rect 53060 54288 53124 54352
rect 53140 54288 53204 54352
rect 53220 54288 53284 54352
rect 58740 54288 58804 54352
rect 58820 54288 58884 54352
rect 58900 54288 58964 54352
rect 58980 54288 59044 54352
rect 59060 54288 59124 54352
rect 59140 54348 59204 54352
rect 59140 54292 59196 54348
rect 59196 54292 59204 54348
rect 59140 54288 59204 54292
rect 59220 54288 59284 54352
rect 64740 54288 64804 54352
rect 64820 54288 64884 54352
rect 64900 54288 64964 54352
rect 64980 54288 65044 54352
rect 65060 54288 65124 54352
rect 65140 54288 65204 54352
rect 65220 54288 65284 54352
rect 70740 54288 70804 54352
rect 70820 54288 70884 54352
rect 70900 54288 70964 54352
rect 70980 54288 71044 54352
rect 71060 54288 71124 54352
rect 71140 54288 71204 54352
rect 71220 54288 71284 54352
rect 1740 52176 1804 52240
rect 1820 52176 1884 52240
rect 1900 52176 1964 52240
rect 1980 52176 2044 52240
rect 2060 52176 2124 52240
rect 2140 52176 2204 52240
rect 2220 52236 2284 52240
rect 2220 52180 2276 52236
rect 2276 52180 2284 52236
rect 2220 52176 2284 52180
rect 7740 52176 7804 52240
rect 7820 52176 7884 52240
rect 7900 52176 7964 52240
rect 7980 52176 8044 52240
rect 8060 52176 8124 52240
rect 8140 52176 8204 52240
rect 8220 52176 8284 52240
rect 13740 52176 13804 52240
rect 13820 52176 13884 52240
rect 13900 52176 13964 52240
rect 13980 52176 14044 52240
rect 14060 52176 14124 52240
rect 14140 52236 14204 52240
rect 14140 52180 14155 52236
rect 14155 52180 14204 52236
rect 14140 52176 14204 52180
rect 14220 52176 14284 52240
rect 19740 52176 19804 52240
rect 19820 52176 19884 52240
rect 19900 52236 19964 52240
rect 19980 52236 20044 52240
rect 19900 52180 19935 52236
rect 19935 52180 19964 52236
rect 19980 52180 19991 52236
rect 19991 52180 20044 52236
rect 19900 52176 19964 52180
rect 19980 52176 20044 52180
rect 20060 52176 20124 52240
rect 20140 52176 20204 52240
rect 20220 52176 20284 52240
rect 25740 52236 25804 52240
rect 25740 52180 25771 52236
rect 25771 52180 25804 52236
rect 25740 52176 25804 52180
rect 25820 52176 25884 52240
rect 25900 52176 25964 52240
rect 25980 52176 26044 52240
rect 26060 52176 26124 52240
rect 26140 52176 26204 52240
rect 26220 52176 26284 52240
rect 31740 52176 31804 52240
rect 31820 52176 31884 52240
rect 31900 52176 31964 52240
rect 31980 52176 32044 52240
rect 32060 52176 32124 52240
rect 32140 52176 32204 52240
rect 32220 52176 32284 52240
rect 37740 52176 37804 52240
rect 37820 52176 37884 52240
rect 37900 52176 37964 52240
rect 37980 52176 38044 52240
rect 38060 52176 38124 52240
rect 38140 52176 38204 52240
rect 38220 52176 38284 52240
rect 43740 52176 43804 52240
rect 43820 52176 43884 52240
rect 43900 52176 43964 52240
rect 43980 52176 44044 52240
rect 44060 52176 44124 52240
rect 44140 52176 44204 52240
rect 44220 52176 44284 52240
rect 49740 52236 49804 52240
rect 49820 52236 49884 52240
rect 49740 52180 49754 52236
rect 49754 52180 49804 52236
rect 49820 52180 49834 52236
rect 49834 52180 49884 52236
rect 49740 52176 49804 52180
rect 49820 52176 49884 52180
rect 49900 52176 49964 52240
rect 49980 52176 50044 52240
rect 50060 52176 50124 52240
rect 50140 52176 50204 52240
rect 50220 52176 50284 52240
rect 55740 52176 55804 52240
rect 55820 52176 55884 52240
rect 55900 52176 55964 52240
rect 55980 52176 56044 52240
rect 56060 52176 56124 52240
rect 56140 52176 56204 52240
rect 56220 52176 56284 52240
rect 61740 52176 61804 52240
rect 61820 52176 61884 52240
rect 61900 52176 61964 52240
rect 61980 52176 62044 52240
rect 62060 52176 62124 52240
rect 62140 52176 62204 52240
rect 62220 52176 62284 52240
rect 67740 52176 67804 52240
rect 67820 52176 67884 52240
rect 67900 52176 67964 52240
rect 67980 52176 68044 52240
rect 68060 52176 68124 52240
rect 68140 52176 68204 52240
rect 68220 52176 68284 52240
rect 73740 52176 73804 52240
rect 73820 52176 73884 52240
rect 73900 52176 73964 52240
rect 73980 52176 74044 52240
rect 74060 52176 74124 52240
rect 74140 52176 74204 52240
rect 74220 52176 74284 52240
rect 1740 52096 1804 52160
rect 1820 52096 1884 52160
rect 1900 52096 1964 52160
rect 1980 52096 2044 52160
rect 2060 52096 2124 52160
rect 2140 52096 2204 52160
rect 2220 52156 2284 52160
rect 2220 52100 2276 52156
rect 2276 52100 2284 52156
rect 2220 52096 2284 52100
rect 7740 52096 7804 52160
rect 7820 52096 7884 52160
rect 7900 52096 7964 52160
rect 7980 52096 8044 52160
rect 8060 52096 8124 52160
rect 8140 52096 8204 52160
rect 8220 52096 8284 52160
rect 13740 52096 13804 52160
rect 13820 52096 13884 52160
rect 13900 52096 13964 52160
rect 13980 52096 14044 52160
rect 14060 52096 14124 52160
rect 14140 52156 14204 52160
rect 14140 52100 14155 52156
rect 14155 52100 14204 52156
rect 14140 52096 14204 52100
rect 14220 52096 14284 52160
rect 19740 52096 19804 52160
rect 19820 52096 19884 52160
rect 19900 52156 19964 52160
rect 19980 52156 20044 52160
rect 19900 52100 19935 52156
rect 19935 52100 19964 52156
rect 19980 52100 19991 52156
rect 19991 52100 20044 52156
rect 19900 52096 19964 52100
rect 19980 52096 20044 52100
rect 20060 52096 20124 52160
rect 20140 52096 20204 52160
rect 20220 52096 20284 52160
rect 25740 52156 25804 52160
rect 25740 52100 25771 52156
rect 25771 52100 25804 52156
rect 25740 52096 25804 52100
rect 25820 52096 25884 52160
rect 25900 52096 25964 52160
rect 25980 52096 26044 52160
rect 26060 52096 26124 52160
rect 26140 52096 26204 52160
rect 26220 52096 26284 52160
rect 31740 52096 31804 52160
rect 31820 52096 31884 52160
rect 31900 52096 31964 52160
rect 31980 52096 32044 52160
rect 32060 52096 32124 52160
rect 32140 52096 32204 52160
rect 32220 52096 32284 52160
rect 37740 52096 37804 52160
rect 37820 52096 37884 52160
rect 37900 52096 37964 52160
rect 37980 52096 38044 52160
rect 38060 52096 38124 52160
rect 38140 52096 38204 52160
rect 38220 52096 38284 52160
rect 43740 52096 43804 52160
rect 43820 52096 43884 52160
rect 43900 52096 43964 52160
rect 43980 52096 44044 52160
rect 44060 52096 44124 52160
rect 44140 52096 44204 52160
rect 44220 52096 44284 52160
rect 49740 52156 49804 52160
rect 49820 52156 49884 52160
rect 49740 52100 49754 52156
rect 49754 52100 49804 52156
rect 49820 52100 49834 52156
rect 49834 52100 49884 52156
rect 49740 52096 49804 52100
rect 49820 52096 49884 52100
rect 49900 52096 49964 52160
rect 49980 52096 50044 52160
rect 50060 52096 50124 52160
rect 50140 52096 50204 52160
rect 50220 52096 50284 52160
rect 55740 52096 55804 52160
rect 55820 52096 55884 52160
rect 55900 52096 55964 52160
rect 55980 52096 56044 52160
rect 56060 52096 56124 52160
rect 56140 52096 56204 52160
rect 56220 52096 56284 52160
rect 61740 52096 61804 52160
rect 61820 52096 61884 52160
rect 61900 52096 61964 52160
rect 61980 52096 62044 52160
rect 62060 52096 62124 52160
rect 62140 52096 62204 52160
rect 62220 52096 62284 52160
rect 67740 52096 67804 52160
rect 67820 52096 67884 52160
rect 67900 52096 67964 52160
rect 67980 52096 68044 52160
rect 68060 52096 68124 52160
rect 68140 52096 68204 52160
rect 68220 52096 68284 52160
rect 73740 52096 73804 52160
rect 73820 52096 73884 52160
rect 73900 52096 73964 52160
rect 73980 52096 74044 52160
rect 74060 52096 74124 52160
rect 74140 52096 74204 52160
rect 74220 52096 74284 52160
rect 1740 52016 1804 52080
rect 1820 52016 1884 52080
rect 1900 52016 1964 52080
rect 1980 52016 2044 52080
rect 2060 52016 2124 52080
rect 2140 52016 2204 52080
rect 2220 52076 2284 52080
rect 2220 52020 2276 52076
rect 2276 52020 2284 52076
rect 2220 52016 2284 52020
rect 7740 52016 7804 52080
rect 7820 52016 7884 52080
rect 7900 52016 7964 52080
rect 7980 52016 8044 52080
rect 8060 52016 8124 52080
rect 8140 52016 8204 52080
rect 8220 52016 8284 52080
rect 13740 52016 13804 52080
rect 13820 52016 13884 52080
rect 13900 52016 13964 52080
rect 13980 52016 14044 52080
rect 14060 52016 14124 52080
rect 14140 52076 14204 52080
rect 14140 52020 14155 52076
rect 14155 52020 14204 52076
rect 14140 52016 14204 52020
rect 14220 52016 14284 52080
rect 19740 52016 19804 52080
rect 19820 52016 19884 52080
rect 19900 52076 19964 52080
rect 19980 52076 20044 52080
rect 19900 52020 19935 52076
rect 19935 52020 19964 52076
rect 19980 52020 19991 52076
rect 19991 52020 20044 52076
rect 19900 52016 19964 52020
rect 19980 52016 20044 52020
rect 20060 52016 20124 52080
rect 20140 52016 20204 52080
rect 20220 52016 20284 52080
rect 25740 52076 25804 52080
rect 25740 52020 25771 52076
rect 25771 52020 25804 52076
rect 25740 52016 25804 52020
rect 25820 52016 25884 52080
rect 25900 52016 25964 52080
rect 25980 52016 26044 52080
rect 26060 52016 26124 52080
rect 26140 52016 26204 52080
rect 26220 52016 26284 52080
rect 31740 52016 31804 52080
rect 31820 52016 31884 52080
rect 31900 52016 31964 52080
rect 31980 52016 32044 52080
rect 32060 52016 32124 52080
rect 32140 52016 32204 52080
rect 32220 52016 32284 52080
rect 37740 52016 37804 52080
rect 37820 52016 37884 52080
rect 37900 52016 37964 52080
rect 37980 52016 38044 52080
rect 38060 52016 38124 52080
rect 38140 52016 38204 52080
rect 38220 52016 38284 52080
rect 43740 52016 43804 52080
rect 43820 52016 43884 52080
rect 43900 52016 43964 52080
rect 43980 52016 44044 52080
rect 44060 52016 44124 52080
rect 44140 52016 44204 52080
rect 44220 52016 44284 52080
rect 49740 52076 49804 52080
rect 49820 52076 49884 52080
rect 49740 52020 49754 52076
rect 49754 52020 49804 52076
rect 49820 52020 49834 52076
rect 49834 52020 49884 52076
rect 49740 52016 49804 52020
rect 49820 52016 49884 52020
rect 49900 52016 49964 52080
rect 49980 52016 50044 52080
rect 50060 52016 50124 52080
rect 50140 52016 50204 52080
rect 50220 52016 50284 52080
rect 55740 52016 55804 52080
rect 55820 52016 55884 52080
rect 55900 52016 55964 52080
rect 55980 52016 56044 52080
rect 56060 52016 56124 52080
rect 56140 52016 56204 52080
rect 56220 52016 56284 52080
rect 61740 52016 61804 52080
rect 61820 52016 61884 52080
rect 61900 52016 61964 52080
rect 61980 52016 62044 52080
rect 62060 52016 62124 52080
rect 62140 52016 62204 52080
rect 62220 52016 62284 52080
rect 67740 52016 67804 52080
rect 67820 52016 67884 52080
rect 67900 52016 67964 52080
rect 67980 52016 68044 52080
rect 68060 52016 68124 52080
rect 68140 52016 68204 52080
rect 68220 52016 68284 52080
rect 73740 52016 73804 52080
rect 73820 52016 73884 52080
rect 73900 52016 73964 52080
rect 73980 52016 74044 52080
rect 74060 52016 74124 52080
rect 74140 52016 74204 52080
rect 74220 52016 74284 52080
rect 1740 51936 1804 52000
rect 1820 51936 1884 52000
rect 1900 51936 1964 52000
rect 1980 51936 2044 52000
rect 2060 51936 2124 52000
rect 2140 51936 2204 52000
rect 2220 51996 2284 52000
rect 2220 51940 2276 51996
rect 2276 51940 2284 51996
rect 2220 51936 2284 51940
rect 7740 51936 7804 52000
rect 7820 51936 7884 52000
rect 7900 51936 7964 52000
rect 7980 51936 8044 52000
rect 8060 51936 8124 52000
rect 8140 51936 8204 52000
rect 8220 51936 8284 52000
rect 13740 51936 13804 52000
rect 13820 51936 13884 52000
rect 13900 51936 13964 52000
rect 13980 51936 14044 52000
rect 14060 51936 14124 52000
rect 14140 51996 14204 52000
rect 14140 51940 14155 51996
rect 14155 51940 14204 51996
rect 14140 51936 14204 51940
rect 14220 51936 14284 52000
rect 19740 51936 19804 52000
rect 19820 51936 19884 52000
rect 19900 51996 19964 52000
rect 19980 51996 20044 52000
rect 19900 51940 19935 51996
rect 19935 51940 19964 51996
rect 19980 51940 19991 51996
rect 19991 51940 20044 51996
rect 19900 51936 19964 51940
rect 19980 51936 20044 51940
rect 20060 51936 20124 52000
rect 20140 51936 20204 52000
rect 20220 51936 20284 52000
rect 25740 51996 25804 52000
rect 25740 51940 25771 51996
rect 25771 51940 25804 51996
rect 25740 51936 25804 51940
rect 25820 51936 25884 52000
rect 25900 51936 25964 52000
rect 25980 51936 26044 52000
rect 26060 51936 26124 52000
rect 26140 51936 26204 52000
rect 26220 51936 26284 52000
rect 31740 51936 31804 52000
rect 31820 51936 31884 52000
rect 31900 51936 31964 52000
rect 31980 51936 32044 52000
rect 32060 51936 32124 52000
rect 32140 51936 32204 52000
rect 32220 51936 32284 52000
rect 37740 51936 37804 52000
rect 37820 51936 37884 52000
rect 37900 51936 37964 52000
rect 37980 51936 38044 52000
rect 38060 51936 38124 52000
rect 38140 51936 38204 52000
rect 38220 51936 38284 52000
rect 43740 51936 43804 52000
rect 43820 51936 43884 52000
rect 43900 51936 43964 52000
rect 43980 51936 44044 52000
rect 44060 51936 44124 52000
rect 44140 51936 44204 52000
rect 44220 51936 44284 52000
rect 49740 51996 49804 52000
rect 49820 51996 49884 52000
rect 49740 51940 49754 51996
rect 49754 51940 49804 51996
rect 49820 51940 49834 51996
rect 49834 51940 49884 51996
rect 49740 51936 49804 51940
rect 49820 51936 49884 51940
rect 49900 51936 49964 52000
rect 49980 51936 50044 52000
rect 50060 51936 50124 52000
rect 50140 51936 50204 52000
rect 50220 51936 50284 52000
rect 55740 51936 55804 52000
rect 55820 51936 55884 52000
rect 55900 51936 55964 52000
rect 55980 51936 56044 52000
rect 56060 51936 56124 52000
rect 56140 51936 56204 52000
rect 56220 51936 56284 52000
rect 61740 51936 61804 52000
rect 61820 51936 61884 52000
rect 61900 51936 61964 52000
rect 61980 51936 62044 52000
rect 62060 51936 62124 52000
rect 62140 51936 62204 52000
rect 62220 51936 62284 52000
rect 67740 51936 67804 52000
rect 67820 51936 67884 52000
rect 67900 51936 67964 52000
rect 67980 51936 68044 52000
rect 68060 51936 68124 52000
rect 68140 51936 68204 52000
rect 68220 51936 68284 52000
rect 73740 51936 73804 52000
rect 73820 51936 73884 52000
rect 73900 51936 73964 52000
rect 73980 51936 74044 52000
rect 74060 51936 74124 52000
rect 74140 51936 74204 52000
rect 74220 51936 74284 52000
rect 65748 47016 65812 47020
rect 65748 46960 65762 47016
rect 65762 46960 65812 47016
rect 65748 46956 65812 46960
rect 66116 46956 66180 47020
rect 4740 44528 4804 44592
rect 4820 44528 4884 44592
rect 4900 44528 4964 44592
rect 4980 44528 5044 44592
rect 5060 44528 5124 44592
rect 5140 44528 5204 44592
rect 5220 44528 5284 44592
rect 10740 44528 10804 44592
rect 10820 44528 10884 44592
rect 10900 44528 10964 44592
rect 10980 44528 11044 44592
rect 11060 44528 11124 44592
rect 11140 44528 11204 44592
rect 11220 44528 11284 44592
rect 16740 44528 16804 44592
rect 16820 44528 16884 44592
rect 16900 44528 16964 44592
rect 16980 44528 17044 44592
rect 17060 44528 17124 44592
rect 17140 44588 17204 44592
rect 17220 44588 17284 44592
rect 17140 44532 17192 44588
rect 17192 44532 17204 44588
rect 17220 44532 17248 44588
rect 17248 44532 17284 44588
rect 17140 44528 17204 44532
rect 17220 44528 17284 44532
rect 22740 44528 22804 44592
rect 22820 44528 22884 44592
rect 22900 44528 22964 44592
rect 22980 44588 23044 44592
rect 22980 44532 23028 44588
rect 23028 44532 23044 44588
rect 22980 44528 23044 44532
rect 23060 44528 23124 44592
rect 23140 44528 23204 44592
rect 23220 44528 23284 44592
rect 28740 44588 28804 44592
rect 28740 44532 28752 44588
rect 28752 44532 28804 44588
rect 28740 44528 28804 44532
rect 28820 44528 28884 44592
rect 28900 44528 28964 44592
rect 28980 44528 29044 44592
rect 29060 44528 29124 44592
rect 29140 44528 29204 44592
rect 29220 44528 29284 44592
rect 34740 44528 34804 44592
rect 34820 44528 34884 44592
rect 34900 44528 34964 44592
rect 34980 44528 35044 44592
rect 35060 44528 35124 44592
rect 35140 44528 35204 44592
rect 35220 44528 35284 44592
rect 40740 44528 40804 44592
rect 40820 44528 40884 44592
rect 40900 44528 40964 44592
rect 40980 44528 41044 44592
rect 41060 44528 41124 44592
rect 41140 44528 41204 44592
rect 41220 44528 41284 44592
rect 46740 44528 46804 44592
rect 46820 44528 46884 44592
rect 46900 44528 46964 44592
rect 46980 44528 47044 44592
rect 47060 44528 47124 44592
rect 47140 44528 47204 44592
rect 47220 44528 47284 44592
rect 52740 44528 52804 44592
rect 52820 44528 52884 44592
rect 52900 44528 52964 44592
rect 52980 44528 53044 44592
rect 53060 44528 53124 44592
rect 53140 44528 53204 44592
rect 53220 44528 53284 44592
rect 58740 44528 58804 44592
rect 58820 44528 58884 44592
rect 58900 44528 58964 44592
rect 58980 44528 59044 44592
rect 59060 44528 59124 44592
rect 59140 44588 59204 44592
rect 59140 44532 59196 44588
rect 59196 44532 59204 44588
rect 59140 44528 59204 44532
rect 59220 44528 59284 44592
rect 64740 44528 64804 44592
rect 64820 44528 64884 44592
rect 64900 44528 64964 44592
rect 64980 44528 65044 44592
rect 65060 44528 65124 44592
rect 65140 44528 65204 44592
rect 65220 44528 65284 44592
rect 70740 44528 70804 44592
rect 70820 44528 70884 44592
rect 70900 44528 70964 44592
rect 70980 44528 71044 44592
rect 71060 44528 71124 44592
rect 71140 44528 71204 44592
rect 71220 44528 71284 44592
rect 4740 44448 4804 44512
rect 4820 44448 4884 44512
rect 4900 44448 4964 44512
rect 4980 44448 5044 44512
rect 5060 44448 5124 44512
rect 5140 44448 5204 44512
rect 5220 44448 5284 44512
rect 10740 44448 10804 44512
rect 10820 44448 10884 44512
rect 10900 44448 10964 44512
rect 10980 44448 11044 44512
rect 11060 44448 11124 44512
rect 11140 44448 11204 44512
rect 11220 44448 11284 44512
rect 16740 44448 16804 44512
rect 16820 44448 16884 44512
rect 16900 44448 16964 44512
rect 16980 44448 17044 44512
rect 17060 44448 17124 44512
rect 17140 44508 17204 44512
rect 17220 44508 17284 44512
rect 17140 44452 17192 44508
rect 17192 44452 17204 44508
rect 17220 44452 17248 44508
rect 17248 44452 17284 44508
rect 17140 44448 17204 44452
rect 17220 44448 17284 44452
rect 22740 44448 22804 44512
rect 22820 44448 22884 44512
rect 22900 44448 22964 44512
rect 22980 44508 23044 44512
rect 22980 44452 23028 44508
rect 23028 44452 23044 44508
rect 22980 44448 23044 44452
rect 23060 44448 23124 44512
rect 23140 44448 23204 44512
rect 23220 44448 23284 44512
rect 28740 44508 28804 44512
rect 28740 44452 28752 44508
rect 28752 44452 28804 44508
rect 28740 44448 28804 44452
rect 28820 44448 28884 44512
rect 28900 44448 28964 44512
rect 28980 44448 29044 44512
rect 29060 44448 29124 44512
rect 29140 44448 29204 44512
rect 29220 44448 29284 44512
rect 34740 44448 34804 44512
rect 34820 44448 34884 44512
rect 34900 44448 34964 44512
rect 34980 44448 35044 44512
rect 35060 44448 35124 44512
rect 35140 44448 35204 44512
rect 35220 44448 35284 44512
rect 40740 44448 40804 44512
rect 40820 44448 40884 44512
rect 40900 44448 40964 44512
rect 40980 44448 41044 44512
rect 41060 44448 41124 44512
rect 41140 44448 41204 44512
rect 41220 44448 41284 44512
rect 46740 44448 46804 44512
rect 46820 44448 46884 44512
rect 46900 44448 46964 44512
rect 46980 44448 47044 44512
rect 47060 44448 47124 44512
rect 47140 44448 47204 44512
rect 47220 44448 47284 44512
rect 52740 44448 52804 44512
rect 52820 44448 52884 44512
rect 52900 44448 52964 44512
rect 52980 44448 53044 44512
rect 53060 44448 53124 44512
rect 53140 44448 53204 44512
rect 53220 44448 53284 44512
rect 58740 44448 58804 44512
rect 58820 44448 58884 44512
rect 58900 44448 58964 44512
rect 58980 44448 59044 44512
rect 59060 44448 59124 44512
rect 59140 44508 59204 44512
rect 59140 44452 59196 44508
rect 59196 44452 59204 44508
rect 59140 44448 59204 44452
rect 59220 44448 59284 44512
rect 64740 44448 64804 44512
rect 64820 44448 64884 44512
rect 64900 44448 64964 44512
rect 64980 44448 65044 44512
rect 65060 44448 65124 44512
rect 65140 44448 65204 44512
rect 65220 44448 65284 44512
rect 70740 44448 70804 44512
rect 70820 44448 70884 44512
rect 70900 44448 70964 44512
rect 70980 44448 71044 44512
rect 71060 44448 71124 44512
rect 71140 44448 71204 44512
rect 71220 44448 71284 44512
rect 4740 44368 4804 44432
rect 4820 44368 4884 44432
rect 4900 44368 4964 44432
rect 4980 44368 5044 44432
rect 5060 44368 5124 44432
rect 5140 44368 5204 44432
rect 5220 44368 5284 44432
rect 10740 44368 10804 44432
rect 10820 44368 10884 44432
rect 10900 44368 10964 44432
rect 10980 44368 11044 44432
rect 11060 44368 11124 44432
rect 11140 44368 11204 44432
rect 11220 44368 11284 44432
rect 16740 44368 16804 44432
rect 16820 44368 16884 44432
rect 16900 44368 16964 44432
rect 16980 44368 17044 44432
rect 17060 44368 17124 44432
rect 17140 44428 17204 44432
rect 17220 44428 17284 44432
rect 17140 44372 17192 44428
rect 17192 44372 17204 44428
rect 17220 44372 17248 44428
rect 17248 44372 17284 44428
rect 17140 44368 17204 44372
rect 17220 44368 17284 44372
rect 22740 44368 22804 44432
rect 22820 44368 22884 44432
rect 22900 44368 22964 44432
rect 22980 44428 23044 44432
rect 22980 44372 23028 44428
rect 23028 44372 23044 44428
rect 22980 44368 23044 44372
rect 23060 44368 23124 44432
rect 23140 44368 23204 44432
rect 23220 44368 23284 44432
rect 28740 44428 28804 44432
rect 28740 44372 28752 44428
rect 28752 44372 28804 44428
rect 28740 44368 28804 44372
rect 28820 44368 28884 44432
rect 28900 44368 28964 44432
rect 28980 44368 29044 44432
rect 29060 44368 29124 44432
rect 29140 44368 29204 44432
rect 29220 44368 29284 44432
rect 34740 44368 34804 44432
rect 34820 44368 34884 44432
rect 34900 44368 34964 44432
rect 34980 44368 35044 44432
rect 35060 44368 35124 44432
rect 35140 44368 35204 44432
rect 35220 44368 35284 44432
rect 40740 44368 40804 44432
rect 40820 44368 40884 44432
rect 40900 44368 40964 44432
rect 40980 44368 41044 44432
rect 41060 44368 41124 44432
rect 41140 44368 41204 44432
rect 41220 44368 41284 44432
rect 46740 44368 46804 44432
rect 46820 44368 46884 44432
rect 46900 44368 46964 44432
rect 46980 44368 47044 44432
rect 47060 44368 47124 44432
rect 47140 44368 47204 44432
rect 47220 44368 47284 44432
rect 52740 44368 52804 44432
rect 52820 44368 52884 44432
rect 52900 44368 52964 44432
rect 52980 44368 53044 44432
rect 53060 44368 53124 44432
rect 53140 44368 53204 44432
rect 53220 44368 53284 44432
rect 58740 44368 58804 44432
rect 58820 44368 58884 44432
rect 58900 44368 58964 44432
rect 58980 44368 59044 44432
rect 59060 44368 59124 44432
rect 59140 44428 59204 44432
rect 59140 44372 59196 44428
rect 59196 44372 59204 44428
rect 59140 44368 59204 44372
rect 59220 44368 59284 44432
rect 64740 44368 64804 44432
rect 64820 44368 64884 44432
rect 64900 44368 64964 44432
rect 64980 44368 65044 44432
rect 65060 44368 65124 44432
rect 65140 44368 65204 44432
rect 65220 44368 65284 44432
rect 70740 44368 70804 44432
rect 70820 44368 70884 44432
rect 70900 44368 70964 44432
rect 70980 44368 71044 44432
rect 71060 44368 71124 44432
rect 71140 44368 71204 44432
rect 71220 44368 71284 44432
rect 4740 44288 4804 44352
rect 4820 44288 4884 44352
rect 4900 44288 4964 44352
rect 4980 44288 5044 44352
rect 5060 44288 5124 44352
rect 5140 44288 5204 44352
rect 5220 44288 5284 44352
rect 10740 44288 10804 44352
rect 10820 44288 10884 44352
rect 10900 44288 10964 44352
rect 10980 44288 11044 44352
rect 11060 44288 11124 44352
rect 11140 44288 11204 44352
rect 11220 44288 11284 44352
rect 16740 44288 16804 44352
rect 16820 44288 16884 44352
rect 16900 44288 16964 44352
rect 16980 44288 17044 44352
rect 17060 44288 17124 44352
rect 17140 44348 17204 44352
rect 17220 44348 17284 44352
rect 17140 44292 17192 44348
rect 17192 44292 17204 44348
rect 17220 44292 17248 44348
rect 17248 44292 17284 44348
rect 17140 44288 17204 44292
rect 17220 44288 17284 44292
rect 22740 44288 22804 44352
rect 22820 44288 22884 44352
rect 22900 44288 22964 44352
rect 22980 44348 23044 44352
rect 22980 44292 23028 44348
rect 23028 44292 23044 44348
rect 22980 44288 23044 44292
rect 23060 44288 23124 44352
rect 23140 44288 23204 44352
rect 23220 44288 23284 44352
rect 28740 44348 28804 44352
rect 28740 44292 28752 44348
rect 28752 44292 28804 44348
rect 28740 44288 28804 44292
rect 28820 44288 28884 44352
rect 28900 44288 28964 44352
rect 28980 44288 29044 44352
rect 29060 44288 29124 44352
rect 29140 44288 29204 44352
rect 29220 44288 29284 44352
rect 34740 44288 34804 44352
rect 34820 44288 34884 44352
rect 34900 44288 34964 44352
rect 34980 44288 35044 44352
rect 35060 44288 35124 44352
rect 35140 44288 35204 44352
rect 35220 44288 35284 44352
rect 40740 44288 40804 44352
rect 40820 44288 40884 44352
rect 40900 44288 40964 44352
rect 40980 44288 41044 44352
rect 41060 44288 41124 44352
rect 41140 44288 41204 44352
rect 41220 44288 41284 44352
rect 46740 44288 46804 44352
rect 46820 44288 46884 44352
rect 46900 44288 46964 44352
rect 46980 44288 47044 44352
rect 47060 44288 47124 44352
rect 47140 44288 47204 44352
rect 47220 44288 47284 44352
rect 52740 44288 52804 44352
rect 52820 44288 52884 44352
rect 52900 44288 52964 44352
rect 52980 44288 53044 44352
rect 53060 44288 53124 44352
rect 53140 44288 53204 44352
rect 53220 44288 53284 44352
rect 58740 44288 58804 44352
rect 58820 44288 58884 44352
rect 58900 44288 58964 44352
rect 58980 44288 59044 44352
rect 59060 44288 59124 44352
rect 59140 44348 59204 44352
rect 59140 44292 59196 44348
rect 59196 44292 59204 44348
rect 59140 44288 59204 44292
rect 59220 44288 59284 44352
rect 64740 44288 64804 44352
rect 64820 44288 64884 44352
rect 64900 44288 64964 44352
rect 64980 44288 65044 44352
rect 65060 44288 65124 44352
rect 65140 44288 65204 44352
rect 65220 44288 65284 44352
rect 70740 44288 70804 44352
rect 70820 44288 70884 44352
rect 70900 44288 70964 44352
rect 70980 44288 71044 44352
rect 71060 44288 71124 44352
rect 71140 44288 71204 44352
rect 71220 44288 71284 44352
rect 1740 42176 1804 42240
rect 1820 42176 1884 42240
rect 1900 42176 1964 42240
rect 1980 42176 2044 42240
rect 2060 42176 2124 42240
rect 2140 42176 2204 42240
rect 2220 42236 2284 42240
rect 2220 42180 2276 42236
rect 2276 42180 2284 42236
rect 2220 42176 2284 42180
rect 7740 42176 7804 42240
rect 7820 42176 7884 42240
rect 7900 42176 7964 42240
rect 7980 42176 8044 42240
rect 8060 42176 8124 42240
rect 8140 42176 8204 42240
rect 8220 42176 8284 42240
rect 13740 42176 13804 42240
rect 13820 42176 13884 42240
rect 13900 42176 13964 42240
rect 13980 42176 14044 42240
rect 14060 42176 14124 42240
rect 14140 42236 14204 42240
rect 14140 42180 14155 42236
rect 14155 42180 14204 42236
rect 14140 42176 14204 42180
rect 14220 42176 14284 42240
rect 19740 42176 19804 42240
rect 19820 42176 19884 42240
rect 19900 42236 19964 42240
rect 19980 42236 20044 42240
rect 19900 42180 19935 42236
rect 19935 42180 19964 42236
rect 19980 42180 19991 42236
rect 19991 42180 20044 42236
rect 19900 42176 19964 42180
rect 19980 42176 20044 42180
rect 20060 42176 20124 42240
rect 20140 42176 20204 42240
rect 20220 42176 20284 42240
rect 25740 42236 25804 42240
rect 25740 42180 25771 42236
rect 25771 42180 25804 42236
rect 25740 42176 25804 42180
rect 25820 42176 25884 42240
rect 25900 42176 25964 42240
rect 25980 42176 26044 42240
rect 26060 42176 26124 42240
rect 26140 42176 26204 42240
rect 26220 42176 26284 42240
rect 31740 42176 31804 42240
rect 31820 42176 31884 42240
rect 31900 42176 31964 42240
rect 31980 42176 32044 42240
rect 32060 42176 32124 42240
rect 32140 42176 32204 42240
rect 32220 42176 32284 42240
rect 37740 42176 37804 42240
rect 37820 42176 37884 42240
rect 37900 42176 37964 42240
rect 37980 42176 38044 42240
rect 38060 42176 38124 42240
rect 38140 42176 38204 42240
rect 38220 42176 38284 42240
rect 43740 42176 43804 42240
rect 43820 42176 43884 42240
rect 43900 42176 43964 42240
rect 43980 42176 44044 42240
rect 44060 42176 44124 42240
rect 44140 42176 44204 42240
rect 44220 42176 44284 42240
rect 49740 42236 49804 42240
rect 49820 42236 49884 42240
rect 49740 42180 49754 42236
rect 49754 42180 49804 42236
rect 49820 42180 49834 42236
rect 49834 42180 49884 42236
rect 49740 42176 49804 42180
rect 49820 42176 49884 42180
rect 49900 42176 49964 42240
rect 49980 42176 50044 42240
rect 50060 42176 50124 42240
rect 50140 42176 50204 42240
rect 50220 42176 50284 42240
rect 55740 42176 55804 42240
rect 55820 42176 55884 42240
rect 55900 42176 55964 42240
rect 55980 42176 56044 42240
rect 56060 42176 56124 42240
rect 56140 42176 56204 42240
rect 56220 42176 56284 42240
rect 61740 42176 61804 42240
rect 61820 42176 61884 42240
rect 61900 42176 61964 42240
rect 61980 42176 62044 42240
rect 62060 42176 62124 42240
rect 62140 42176 62204 42240
rect 62220 42176 62284 42240
rect 67740 42176 67804 42240
rect 67820 42176 67884 42240
rect 67900 42176 67964 42240
rect 67980 42176 68044 42240
rect 68060 42176 68124 42240
rect 68140 42176 68204 42240
rect 68220 42176 68284 42240
rect 73740 42176 73804 42240
rect 73820 42176 73884 42240
rect 73900 42176 73964 42240
rect 73980 42176 74044 42240
rect 74060 42176 74124 42240
rect 74140 42176 74204 42240
rect 74220 42176 74284 42240
rect 1740 42096 1804 42160
rect 1820 42096 1884 42160
rect 1900 42096 1964 42160
rect 1980 42096 2044 42160
rect 2060 42096 2124 42160
rect 2140 42096 2204 42160
rect 2220 42156 2284 42160
rect 2220 42100 2276 42156
rect 2276 42100 2284 42156
rect 2220 42096 2284 42100
rect 7740 42096 7804 42160
rect 7820 42096 7884 42160
rect 7900 42096 7964 42160
rect 7980 42096 8044 42160
rect 8060 42096 8124 42160
rect 8140 42096 8204 42160
rect 8220 42096 8284 42160
rect 13740 42096 13804 42160
rect 13820 42096 13884 42160
rect 13900 42096 13964 42160
rect 13980 42096 14044 42160
rect 14060 42096 14124 42160
rect 14140 42156 14204 42160
rect 14140 42100 14155 42156
rect 14155 42100 14204 42156
rect 14140 42096 14204 42100
rect 14220 42096 14284 42160
rect 19740 42096 19804 42160
rect 19820 42096 19884 42160
rect 19900 42156 19964 42160
rect 19980 42156 20044 42160
rect 19900 42100 19935 42156
rect 19935 42100 19964 42156
rect 19980 42100 19991 42156
rect 19991 42100 20044 42156
rect 19900 42096 19964 42100
rect 19980 42096 20044 42100
rect 20060 42096 20124 42160
rect 20140 42096 20204 42160
rect 20220 42096 20284 42160
rect 25740 42156 25804 42160
rect 25740 42100 25771 42156
rect 25771 42100 25804 42156
rect 25740 42096 25804 42100
rect 25820 42096 25884 42160
rect 25900 42096 25964 42160
rect 25980 42096 26044 42160
rect 26060 42096 26124 42160
rect 26140 42096 26204 42160
rect 26220 42096 26284 42160
rect 31740 42096 31804 42160
rect 31820 42096 31884 42160
rect 31900 42096 31964 42160
rect 31980 42096 32044 42160
rect 32060 42096 32124 42160
rect 32140 42096 32204 42160
rect 32220 42096 32284 42160
rect 37740 42096 37804 42160
rect 37820 42096 37884 42160
rect 37900 42096 37964 42160
rect 37980 42096 38044 42160
rect 38060 42096 38124 42160
rect 38140 42096 38204 42160
rect 38220 42096 38284 42160
rect 43740 42096 43804 42160
rect 43820 42096 43884 42160
rect 43900 42096 43964 42160
rect 43980 42096 44044 42160
rect 44060 42096 44124 42160
rect 44140 42096 44204 42160
rect 44220 42096 44284 42160
rect 49740 42156 49804 42160
rect 49820 42156 49884 42160
rect 49740 42100 49754 42156
rect 49754 42100 49804 42156
rect 49820 42100 49834 42156
rect 49834 42100 49884 42156
rect 49740 42096 49804 42100
rect 49820 42096 49884 42100
rect 49900 42096 49964 42160
rect 49980 42096 50044 42160
rect 50060 42096 50124 42160
rect 50140 42096 50204 42160
rect 50220 42096 50284 42160
rect 55740 42096 55804 42160
rect 55820 42096 55884 42160
rect 55900 42096 55964 42160
rect 55980 42096 56044 42160
rect 56060 42096 56124 42160
rect 56140 42096 56204 42160
rect 56220 42096 56284 42160
rect 61740 42096 61804 42160
rect 61820 42096 61884 42160
rect 61900 42096 61964 42160
rect 61980 42096 62044 42160
rect 62060 42096 62124 42160
rect 62140 42096 62204 42160
rect 62220 42096 62284 42160
rect 67740 42096 67804 42160
rect 67820 42096 67884 42160
rect 67900 42096 67964 42160
rect 67980 42096 68044 42160
rect 68060 42096 68124 42160
rect 68140 42096 68204 42160
rect 68220 42096 68284 42160
rect 73740 42096 73804 42160
rect 73820 42096 73884 42160
rect 73900 42096 73964 42160
rect 73980 42096 74044 42160
rect 74060 42096 74124 42160
rect 74140 42096 74204 42160
rect 74220 42096 74284 42160
rect 1740 42016 1804 42080
rect 1820 42016 1884 42080
rect 1900 42016 1964 42080
rect 1980 42016 2044 42080
rect 2060 42016 2124 42080
rect 2140 42016 2204 42080
rect 2220 42076 2284 42080
rect 2220 42020 2276 42076
rect 2276 42020 2284 42076
rect 2220 42016 2284 42020
rect 7740 42016 7804 42080
rect 7820 42016 7884 42080
rect 7900 42016 7964 42080
rect 7980 42016 8044 42080
rect 8060 42016 8124 42080
rect 8140 42016 8204 42080
rect 8220 42016 8284 42080
rect 13740 42016 13804 42080
rect 13820 42016 13884 42080
rect 13900 42016 13964 42080
rect 13980 42016 14044 42080
rect 14060 42016 14124 42080
rect 14140 42076 14204 42080
rect 14140 42020 14155 42076
rect 14155 42020 14204 42076
rect 14140 42016 14204 42020
rect 14220 42016 14284 42080
rect 19740 42016 19804 42080
rect 19820 42016 19884 42080
rect 19900 42076 19964 42080
rect 19980 42076 20044 42080
rect 19900 42020 19935 42076
rect 19935 42020 19964 42076
rect 19980 42020 19991 42076
rect 19991 42020 20044 42076
rect 19900 42016 19964 42020
rect 19980 42016 20044 42020
rect 20060 42016 20124 42080
rect 20140 42016 20204 42080
rect 20220 42016 20284 42080
rect 25740 42076 25804 42080
rect 25740 42020 25771 42076
rect 25771 42020 25804 42076
rect 25740 42016 25804 42020
rect 25820 42016 25884 42080
rect 25900 42016 25964 42080
rect 25980 42016 26044 42080
rect 26060 42016 26124 42080
rect 26140 42016 26204 42080
rect 26220 42016 26284 42080
rect 31740 42016 31804 42080
rect 31820 42016 31884 42080
rect 31900 42016 31964 42080
rect 31980 42016 32044 42080
rect 32060 42016 32124 42080
rect 32140 42016 32204 42080
rect 32220 42016 32284 42080
rect 37740 42016 37804 42080
rect 37820 42016 37884 42080
rect 37900 42016 37964 42080
rect 37980 42016 38044 42080
rect 38060 42016 38124 42080
rect 38140 42016 38204 42080
rect 38220 42016 38284 42080
rect 43740 42016 43804 42080
rect 43820 42016 43884 42080
rect 43900 42016 43964 42080
rect 43980 42016 44044 42080
rect 44060 42016 44124 42080
rect 44140 42016 44204 42080
rect 44220 42016 44284 42080
rect 49740 42076 49804 42080
rect 49820 42076 49884 42080
rect 49740 42020 49754 42076
rect 49754 42020 49804 42076
rect 49820 42020 49834 42076
rect 49834 42020 49884 42076
rect 49740 42016 49804 42020
rect 49820 42016 49884 42020
rect 49900 42016 49964 42080
rect 49980 42016 50044 42080
rect 50060 42016 50124 42080
rect 50140 42016 50204 42080
rect 50220 42016 50284 42080
rect 55740 42016 55804 42080
rect 55820 42016 55884 42080
rect 55900 42016 55964 42080
rect 55980 42016 56044 42080
rect 56060 42016 56124 42080
rect 56140 42016 56204 42080
rect 56220 42016 56284 42080
rect 61740 42016 61804 42080
rect 61820 42016 61884 42080
rect 61900 42016 61964 42080
rect 61980 42016 62044 42080
rect 62060 42016 62124 42080
rect 62140 42016 62204 42080
rect 62220 42016 62284 42080
rect 67740 42016 67804 42080
rect 67820 42016 67884 42080
rect 67900 42016 67964 42080
rect 67980 42016 68044 42080
rect 68060 42016 68124 42080
rect 68140 42016 68204 42080
rect 68220 42016 68284 42080
rect 73740 42016 73804 42080
rect 73820 42016 73884 42080
rect 73900 42016 73964 42080
rect 73980 42016 74044 42080
rect 74060 42016 74124 42080
rect 74140 42016 74204 42080
rect 74220 42016 74284 42080
rect 1740 41936 1804 42000
rect 1820 41936 1884 42000
rect 1900 41936 1964 42000
rect 1980 41936 2044 42000
rect 2060 41936 2124 42000
rect 2140 41936 2204 42000
rect 2220 41996 2284 42000
rect 2220 41940 2276 41996
rect 2276 41940 2284 41996
rect 2220 41936 2284 41940
rect 7740 41936 7804 42000
rect 7820 41936 7884 42000
rect 7900 41936 7964 42000
rect 7980 41936 8044 42000
rect 8060 41936 8124 42000
rect 8140 41936 8204 42000
rect 8220 41936 8284 42000
rect 13740 41936 13804 42000
rect 13820 41936 13884 42000
rect 13900 41936 13964 42000
rect 13980 41936 14044 42000
rect 14060 41936 14124 42000
rect 14140 41996 14204 42000
rect 14140 41940 14155 41996
rect 14155 41940 14204 41996
rect 14140 41936 14204 41940
rect 14220 41936 14284 42000
rect 19740 41936 19804 42000
rect 19820 41936 19884 42000
rect 19900 41996 19964 42000
rect 19980 41996 20044 42000
rect 19900 41940 19935 41996
rect 19935 41940 19964 41996
rect 19980 41940 19991 41996
rect 19991 41940 20044 41996
rect 19900 41936 19964 41940
rect 19980 41936 20044 41940
rect 20060 41936 20124 42000
rect 20140 41936 20204 42000
rect 20220 41936 20284 42000
rect 25740 41996 25804 42000
rect 25740 41940 25771 41996
rect 25771 41940 25804 41996
rect 25740 41936 25804 41940
rect 25820 41936 25884 42000
rect 25900 41936 25964 42000
rect 25980 41936 26044 42000
rect 26060 41936 26124 42000
rect 26140 41936 26204 42000
rect 26220 41936 26284 42000
rect 31740 41936 31804 42000
rect 31820 41936 31884 42000
rect 31900 41936 31964 42000
rect 31980 41936 32044 42000
rect 32060 41936 32124 42000
rect 32140 41936 32204 42000
rect 32220 41936 32284 42000
rect 37740 41936 37804 42000
rect 37820 41936 37884 42000
rect 37900 41936 37964 42000
rect 37980 41936 38044 42000
rect 38060 41936 38124 42000
rect 38140 41936 38204 42000
rect 38220 41936 38284 42000
rect 43740 41936 43804 42000
rect 43820 41936 43884 42000
rect 43900 41936 43964 42000
rect 43980 41936 44044 42000
rect 44060 41936 44124 42000
rect 44140 41936 44204 42000
rect 44220 41936 44284 42000
rect 49740 41996 49804 42000
rect 49820 41996 49884 42000
rect 49740 41940 49754 41996
rect 49754 41940 49804 41996
rect 49820 41940 49834 41996
rect 49834 41940 49884 41996
rect 49740 41936 49804 41940
rect 49820 41936 49884 41940
rect 49900 41936 49964 42000
rect 49980 41936 50044 42000
rect 50060 41936 50124 42000
rect 50140 41936 50204 42000
rect 50220 41936 50284 42000
rect 55740 41936 55804 42000
rect 55820 41936 55884 42000
rect 55900 41936 55964 42000
rect 55980 41936 56044 42000
rect 56060 41936 56124 42000
rect 56140 41936 56204 42000
rect 56220 41936 56284 42000
rect 61740 41936 61804 42000
rect 61820 41936 61884 42000
rect 61900 41936 61964 42000
rect 61980 41936 62044 42000
rect 62060 41936 62124 42000
rect 62140 41936 62204 42000
rect 62220 41936 62284 42000
rect 67740 41936 67804 42000
rect 67820 41936 67884 42000
rect 67900 41936 67964 42000
rect 67980 41936 68044 42000
rect 68060 41936 68124 42000
rect 68140 41936 68204 42000
rect 68220 41936 68284 42000
rect 73740 41936 73804 42000
rect 73820 41936 73884 42000
rect 73900 41936 73964 42000
rect 73980 41936 74044 42000
rect 74060 41936 74124 42000
rect 74140 41936 74204 42000
rect 74220 41936 74284 42000
rect 65564 41244 65628 41308
rect 65564 38524 65628 38588
rect 65564 34716 65628 34780
rect 4740 34528 4804 34592
rect 4820 34528 4884 34592
rect 4900 34528 4964 34592
rect 4980 34528 5044 34592
rect 5060 34528 5124 34592
rect 5140 34528 5204 34592
rect 5220 34528 5284 34592
rect 10740 34528 10804 34592
rect 10820 34528 10884 34592
rect 10900 34528 10964 34592
rect 10980 34528 11044 34592
rect 11060 34528 11124 34592
rect 11140 34528 11204 34592
rect 11220 34528 11284 34592
rect 16740 34528 16804 34592
rect 16820 34528 16884 34592
rect 16900 34528 16964 34592
rect 16980 34528 17044 34592
rect 17060 34528 17124 34592
rect 17140 34588 17204 34592
rect 17220 34588 17284 34592
rect 17140 34532 17192 34588
rect 17192 34532 17204 34588
rect 17220 34532 17248 34588
rect 17248 34532 17284 34588
rect 17140 34528 17204 34532
rect 17220 34528 17284 34532
rect 22740 34528 22804 34592
rect 22820 34528 22884 34592
rect 22900 34528 22964 34592
rect 22980 34588 23044 34592
rect 22980 34532 23028 34588
rect 23028 34532 23044 34588
rect 22980 34528 23044 34532
rect 23060 34528 23124 34592
rect 23140 34528 23204 34592
rect 23220 34528 23284 34592
rect 28740 34588 28804 34592
rect 28740 34532 28752 34588
rect 28752 34532 28804 34588
rect 28740 34528 28804 34532
rect 28820 34528 28884 34592
rect 28900 34528 28964 34592
rect 28980 34528 29044 34592
rect 29060 34528 29124 34592
rect 29140 34528 29204 34592
rect 29220 34528 29284 34592
rect 34740 34528 34804 34592
rect 34820 34528 34884 34592
rect 34900 34528 34964 34592
rect 34980 34528 35044 34592
rect 35060 34528 35124 34592
rect 35140 34528 35204 34592
rect 35220 34528 35284 34592
rect 40740 34528 40804 34592
rect 40820 34528 40884 34592
rect 40900 34528 40964 34592
rect 40980 34528 41044 34592
rect 41060 34528 41124 34592
rect 41140 34528 41204 34592
rect 41220 34528 41284 34592
rect 46740 34528 46804 34592
rect 46820 34528 46884 34592
rect 46900 34528 46964 34592
rect 46980 34528 47044 34592
rect 47060 34528 47124 34592
rect 47140 34528 47204 34592
rect 47220 34528 47284 34592
rect 52740 34528 52804 34592
rect 52820 34528 52884 34592
rect 52900 34528 52964 34592
rect 52980 34528 53044 34592
rect 53060 34528 53124 34592
rect 53140 34528 53204 34592
rect 53220 34528 53284 34592
rect 58740 34528 58804 34592
rect 58820 34528 58884 34592
rect 58900 34528 58964 34592
rect 58980 34528 59044 34592
rect 59060 34528 59124 34592
rect 59140 34588 59204 34592
rect 59140 34532 59196 34588
rect 59196 34532 59204 34588
rect 59140 34528 59204 34532
rect 59220 34528 59284 34592
rect 64740 34528 64804 34592
rect 64820 34528 64884 34592
rect 64900 34528 64964 34592
rect 64980 34528 65044 34592
rect 65060 34528 65124 34592
rect 65140 34528 65204 34592
rect 65220 34528 65284 34592
rect 70740 34528 70804 34592
rect 70820 34528 70884 34592
rect 70900 34528 70964 34592
rect 70980 34528 71044 34592
rect 71060 34528 71124 34592
rect 71140 34528 71204 34592
rect 71220 34528 71284 34592
rect 4740 34448 4804 34512
rect 4820 34448 4884 34512
rect 4900 34448 4964 34512
rect 4980 34448 5044 34512
rect 5060 34448 5124 34512
rect 5140 34448 5204 34512
rect 5220 34448 5284 34512
rect 10740 34448 10804 34512
rect 10820 34448 10884 34512
rect 10900 34448 10964 34512
rect 10980 34448 11044 34512
rect 11060 34448 11124 34512
rect 11140 34448 11204 34512
rect 11220 34448 11284 34512
rect 16740 34448 16804 34512
rect 16820 34448 16884 34512
rect 16900 34448 16964 34512
rect 16980 34448 17044 34512
rect 17060 34448 17124 34512
rect 17140 34508 17204 34512
rect 17220 34508 17284 34512
rect 17140 34452 17192 34508
rect 17192 34452 17204 34508
rect 17220 34452 17248 34508
rect 17248 34452 17284 34508
rect 17140 34448 17204 34452
rect 17220 34448 17284 34452
rect 22740 34448 22804 34512
rect 22820 34448 22884 34512
rect 22900 34448 22964 34512
rect 22980 34508 23044 34512
rect 22980 34452 23028 34508
rect 23028 34452 23044 34508
rect 22980 34448 23044 34452
rect 23060 34448 23124 34512
rect 23140 34448 23204 34512
rect 23220 34448 23284 34512
rect 28740 34508 28804 34512
rect 28740 34452 28752 34508
rect 28752 34452 28804 34508
rect 28740 34448 28804 34452
rect 28820 34448 28884 34512
rect 28900 34448 28964 34512
rect 28980 34448 29044 34512
rect 29060 34448 29124 34512
rect 29140 34448 29204 34512
rect 29220 34448 29284 34512
rect 34740 34448 34804 34512
rect 34820 34448 34884 34512
rect 34900 34448 34964 34512
rect 34980 34448 35044 34512
rect 35060 34448 35124 34512
rect 35140 34448 35204 34512
rect 35220 34448 35284 34512
rect 40740 34448 40804 34512
rect 40820 34448 40884 34512
rect 40900 34448 40964 34512
rect 40980 34448 41044 34512
rect 41060 34448 41124 34512
rect 41140 34448 41204 34512
rect 41220 34448 41284 34512
rect 46740 34448 46804 34512
rect 46820 34448 46884 34512
rect 46900 34448 46964 34512
rect 46980 34448 47044 34512
rect 47060 34448 47124 34512
rect 47140 34448 47204 34512
rect 47220 34448 47284 34512
rect 52740 34448 52804 34512
rect 52820 34448 52884 34512
rect 52900 34448 52964 34512
rect 52980 34448 53044 34512
rect 53060 34448 53124 34512
rect 53140 34448 53204 34512
rect 53220 34448 53284 34512
rect 58740 34448 58804 34512
rect 58820 34448 58884 34512
rect 58900 34448 58964 34512
rect 58980 34448 59044 34512
rect 59060 34448 59124 34512
rect 59140 34508 59204 34512
rect 59140 34452 59196 34508
rect 59196 34452 59204 34508
rect 59140 34448 59204 34452
rect 59220 34448 59284 34512
rect 64740 34448 64804 34512
rect 64820 34448 64884 34512
rect 64900 34448 64964 34512
rect 64980 34448 65044 34512
rect 65060 34448 65124 34512
rect 65140 34448 65204 34512
rect 65220 34448 65284 34512
rect 70740 34448 70804 34512
rect 70820 34448 70884 34512
rect 70900 34448 70964 34512
rect 70980 34448 71044 34512
rect 71060 34448 71124 34512
rect 71140 34448 71204 34512
rect 71220 34448 71284 34512
rect 4740 34368 4804 34432
rect 4820 34368 4884 34432
rect 4900 34368 4964 34432
rect 4980 34368 5044 34432
rect 5060 34368 5124 34432
rect 5140 34368 5204 34432
rect 5220 34368 5284 34432
rect 10740 34368 10804 34432
rect 10820 34368 10884 34432
rect 10900 34368 10964 34432
rect 10980 34368 11044 34432
rect 11060 34368 11124 34432
rect 11140 34368 11204 34432
rect 11220 34368 11284 34432
rect 16740 34368 16804 34432
rect 16820 34368 16884 34432
rect 16900 34368 16964 34432
rect 16980 34368 17044 34432
rect 17060 34368 17124 34432
rect 17140 34428 17204 34432
rect 17220 34428 17284 34432
rect 17140 34372 17192 34428
rect 17192 34372 17204 34428
rect 17220 34372 17248 34428
rect 17248 34372 17284 34428
rect 17140 34368 17204 34372
rect 17220 34368 17284 34372
rect 22740 34368 22804 34432
rect 22820 34368 22884 34432
rect 22900 34368 22964 34432
rect 22980 34428 23044 34432
rect 22980 34372 23028 34428
rect 23028 34372 23044 34428
rect 22980 34368 23044 34372
rect 23060 34368 23124 34432
rect 23140 34368 23204 34432
rect 23220 34368 23284 34432
rect 28740 34428 28804 34432
rect 28740 34372 28752 34428
rect 28752 34372 28804 34428
rect 28740 34368 28804 34372
rect 28820 34368 28884 34432
rect 28900 34368 28964 34432
rect 28980 34368 29044 34432
rect 29060 34368 29124 34432
rect 29140 34368 29204 34432
rect 29220 34368 29284 34432
rect 34740 34368 34804 34432
rect 34820 34368 34884 34432
rect 34900 34368 34964 34432
rect 34980 34368 35044 34432
rect 35060 34368 35124 34432
rect 35140 34368 35204 34432
rect 35220 34368 35284 34432
rect 40740 34368 40804 34432
rect 40820 34368 40884 34432
rect 40900 34368 40964 34432
rect 40980 34368 41044 34432
rect 41060 34368 41124 34432
rect 41140 34368 41204 34432
rect 41220 34368 41284 34432
rect 46740 34368 46804 34432
rect 46820 34368 46884 34432
rect 46900 34368 46964 34432
rect 46980 34368 47044 34432
rect 47060 34368 47124 34432
rect 47140 34368 47204 34432
rect 47220 34368 47284 34432
rect 52740 34368 52804 34432
rect 52820 34368 52884 34432
rect 52900 34368 52964 34432
rect 52980 34368 53044 34432
rect 53060 34368 53124 34432
rect 53140 34368 53204 34432
rect 53220 34368 53284 34432
rect 58740 34368 58804 34432
rect 58820 34368 58884 34432
rect 58900 34368 58964 34432
rect 58980 34368 59044 34432
rect 59060 34368 59124 34432
rect 59140 34428 59204 34432
rect 59140 34372 59196 34428
rect 59196 34372 59204 34428
rect 59140 34368 59204 34372
rect 59220 34368 59284 34432
rect 64740 34368 64804 34432
rect 64820 34368 64884 34432
rect 64900 34368 64964 34432
rect 64980 34368 65044 34432
rect 65060 34368 65124 34432
rect 65140 34368 65204 34432
rect 65220 34368 65284 34432
rect 70740 34368 70804 34432
rect 70820 34368 70884 34432
rect 70900 34368 70964 34432
rect 70980 34368 71044 34432
rect 71060 34368 71124 34432
rect 71140 34368 71204 34432
rect 71220 34368 71284 34432
rect 4740 34288 4804 34352
rect 4820 34288 4884 34352
rect 4900 34288 4964 34352
rect 4980 34288 5044 34352
rect 5060 34288 5124 34352
rect 5140 34288 5204 34352
rect 5220 34288 5284 34352
rect 10740 34288 10804 34352
rect 10820 34288 10884 34352
rect 10900 34288 10964 34352
rect 10980 34288 11044 34352
rect 11060 34288 11124 34352
rect 11140 34288 11204 34352
rect 11220 34288 11284 34352
rect 16740 34288 16804 34352
rect 16820 34288 16884 34352
rect 16900 34288 16964 34352
rect 16980 34288 17044 34352
rect 17060 34288 17124 34352
rect 17140 34348 17204 34352
rect 17220 34348 17284 34352
rect 17140 34292 17192 34348
rect 17192 34292 17204 34348
rect 17220 34292 17248 34348
rect 17248 34292 17284 34348
rect 17140 34288 17204 34292
rect 17220 34288 17284 34292
rect 22740 34288 22804 34352
rect 22820 34288 22884 34352
rect 22900 34288 22964 34352
rect 22980 34348 23044 34352
rect 22980 34292 23028 34348
rect 23028 34292 23044 34348
rect 22980 34288 23044 34292
rect 23060 34288 23124 34352
rect 23140 34288 23204 34352
rect 23220 34288 23284 34352
rect 28740 34348 28804 34352
rect 28740 34292 28752 34348
rect 28752 34292 28804 34348
rect 28740 34288 28804 34292
rect 28820 34288 28884 34352
rect 28900 34288 28964 34352
rect 28980 34288 29044 34352
rect 29060 34288 29124 34352
rect 29140 34288 29204 34352
rect 29220 34288 29284 34352
rect 34740 34288 34804 34352
rect 34820 34288 34884 34352
rect 34900 34288 34964 34352
rect 34980 34288 35044 34352
rect 35060 34288 35124 34352
rect 35140 34288 35204 34352
rect 35220 34288 35284 34352
rect 40740 34288 40804 34352
rect 40820 34288 40884 34352
rect 40900 34288 40964 34352
rect 40980 34288 41044 34352
rect 41060 34288 41124 34352
rect 41140 34288 41204 34352
rect 41220 34288 41284 34352
rect 46740 34288 46804 34352
rect 46820 34288 46884 34352
rect 46900 34288 46964 34352
rect 46980 34288 47044 34352
rect 47060 34288 47124 34352
rect 47140 34288 47204 34352
rect 47220 34288 47284 34352
rect 52740 34288 52804 34352
rect 52820 34288 52884 34352
rect 52900 34288 52964 34352
rect 52980 34288 53044 34352
rect 53060 34288 53124 34352
rect 53140 34288 53204 34352
rect 53220 34288 53284 34352
rect 58740 34288 58804 34352
rect 58820 34288 58884 34352
rect 58900 34288 58964 34352
rect 58980 34288 59044 34352
rect 59060 34288 59124 34352
rect 59140 34348 59204 34352
rect 59140 34292 59196 34348
rect 59196 34292 59204 34348
rect 59140 34288 59204 34292
rect 59220 34288 59284 34352
rect 64740 34288 64804 34352
rect 64820 34288 64884 34352
rect 64900 34288 64964 34352
rect 64980 34288 65044 34352
rect 65060 34288 65124 34352
rect 65140 34288 65204 34352
rect 65220 34288 65284 34352
rect 70740 34288 70804 34352
rect 70820 34288 70884 34352
rect 70900 34288 70964 34352
rect 70980 34288 71044 34352
rect 71060 34288 71124 34352
rect 71140 34288 71204 34352
rect 71220 34288 71284 34352
rect 1740 32176 1804 32240
rect 1820 32176 1884 32240
rect 1900 32176 1964 32240
rect 1980 32176 2044 32240
rect 2060 32176 2124 32240
rect 2140 32176 2204 32240
rect 2220 32236 2284 32240
rect 2220 32180 2276 32236
rect 2276 32180 2284 32236
rect 2220 32176 2284 32180
rect 7740 32176 7804 32240
rect 7820 32176 7884 32240
rect 7900 32176 7964 32240
rect 7980 32176 8044 32240
rect 8060 32176 8124 32240
rect 8140 32176 8204 32240
rect 8220 32176 8284 32240
rect 13740 32176 13804 32240
rect 13820 32176 13884 32240
rect 13900 32176 13964 32240
rect 13980 32176 14044 32240
rect 14060 32176 14124 32240
rect 14140 32236 14204 32240
rect 14140 32180 14155 32236
rect 14155 32180 14204 32236
rect 14140 32176 14204 32180
rect 14220 32176 14284 32240
rect 19740 32176 19804 32240
rect 19820 32176 19884 32240
rect 19900 32236 19964 32240
rect 19980 32236 20044 32240
rect 19900 32180 19935 32236
rect 19935 32180 19964 32236
rect 19980 32180 19991 32236
rect 19991 32180 20044 32236
rect 19900 32176 19964 32180
rect 19980 32176 20044 32180
rect 20060 32176 20124 32240
rect 20140 32176 20204 32240
rect 20220 32176 20284 32240
rect 25740 32236 25804 32240
rect 25740 32180 25771 32236
rect 25771 32180 25804 32236
rect 25740 32176 25804 32180
rect 25820 32176 25884 32240
rect 25900 32176 25964 32240
rect 25980 32176 26044 32240
rect 26060 32176 26124 32240
rect 26140 32176 26204 32240
rect 26220 32176 26284 32240
rect 31740 32176 31804 32240
rect 31820 32176 31884 32240
rect 31900 32176 31964 32240
rect 31980 32176 32044 32240
rect 32060 32176 32124 32240
rect 32140 32176 32204 32240
rect 32220 32176 32284 32240
rect 37740 32176 37804 32240
rect 37820 32176 37884 32240
rect 37900 32176 37964 32240
rect 37980 32176 38044 32240
rect 38060 32176 38124 32240
rect 38140 32176 38204 32240
rect 38220 32176 38284 32240
rect 43740 32176 43804 32240
rect 43820 32176 43884 32240
rect 43900 32176 43964 32240
rect 43980 32176 44044 32240
rect 44060 32176 44124 32240
rect 44140 32176 44204 32240
rect 44220 32176 44284 32240
rect 49740 32236 49804 32240
rect 49820 32236 49884 32240
rect 49740 32180 49754 32236
rect 49754 32180 49804 32236
rect 49820 32180 49834 32236
rect 49834 32180 49884 32236
rect 49740 32176 49804 32180
rect 49820 32176 49884 32180
rect 49900 32176 49964 32240
rect 49980 32176 50044 32240
rect 50060 32176 50124 32240
rect 50140 32176 50204 32240
rect 50220 32176 50284 32240
rect 55740 32176 55804 32240
rect 55820 32176 55884 32240
rect 55900 32176 55964 32240
rect 55980 32176 56044 32240
rect 56060 32176 56124 32240
rect 56140 32176 56204 32240
rect 56220 32176 56284 32240
rect 61740 32176 61804 32240
rect 61820 32176 61884 32240
rect 61900 32176 61964 32240
rect 61980 32176 62044 32240
rect 62060 32176 62124 32240
rect 62140 32176 62204 32240
rect 62220 32176 62284 32240
rect 67740 32176 67804 32240
rect 67820 32176 67884 32240
rect 67900 32176 67964 32240
rect 67980 32176 68044 32240
rect 68060 32176 68124 32240
rect 68140 32176 68204 32240
rect 68220 32176 68284 32240
rect 73740 32176 73804 32240
rect 73820 32176 73884 32240
rect 73900 32176 73964 32240
rect 73980 32176 74044 32240
rect 74060 32176 74124 32240
rect 74140 32176 74204 32240
rect 74220 32176 74284 32240
rect 1740 32096 1804 32160
rect 1820 32096 1884 32160
rect 1900 32096 1964 32160
rect 1980 32096 2044 32160
rect 2060 32096 2124 32160
rect 2140 32096 2204 32160
rect 2220 32156 2284 32160
rect 2220 32100 2276 32156
rect 2276 32100 2284 32156
rect 2220 32096 2284 32100
rect 7740 32096 7804 32160
rect 7820 32096 7884 32160
rect 7900 32096 7964 32160
rect 7980 32096 8044 32160
rect 8060 32096 8124 32160
rect 8140 32096 8204 32160
rect 8220 32096 8284 32160
rect 13740 32096 13804 32160
rect 13820 32096 13884 32160
rect 13900 32096 13964 32160
rect 13980 32096 14044 32160
rect 14060 32096 14124 32160
rect 14140 32156 14204 32160
rect 14140 32100 14155 32156
rect 14155 32100 14204 32156
rect 14140 32096 14204 32100
rect 14220 32096 14284 32160
rect 19740 32096 19804 32160
rect 19820 32096 19884 32160
rect 19900 32156 19964 32160
rect 19980 32156 20044 32160
rect 19900 32100 19935 32156
rect 19935 32100 19964 32156
rect 19980 32100 19991 32156
rect 19991 32100 20044 32156
rect 19900 32096 19964 32100
rect 19980 32096 20044 32100
rect 20060 32096 20124 32160
rect 20140 32096 20204 32160
rect 20220 32096 20284 32160
rect 25740 32156 25804 32160
rect 25740 32100 25771 32156
rect 25771 32100 25804 32156
rect 25740 32096 25804 32100
rect 25820 32096 25884 32160
rect 25900 32096 25964 32160
rect 25980 32096 26044 32160
rect 26060 32096 26124 32160
rect 26140 32096 26204 32160
rect 26220 32096 26284 32160
rect 31740 32096 31804 32160
rect 31820 32096 31884 32160
rect 31900 32096 31964 32160
rect 31980 32096 32044 32160
rect 32060 32096 32124 32160
rect 32140 32096 32204 32160
rect 32220 32096 32284 32160
rect 37740 32096 37804 32160
rect 37820 32096 37884 32160
rect 37900 32096 37964 32160
rect 37980 32096 38044 32160
rect 38060 32096 38124 32160
rect 38140 32096 38204 32160
rect 38220 32096 38284 32160
rect 43740 32096 43804 32160
rect 43820 32096 43884 32160
rect 43900 32096 43964 32160
rect 43980 32096 44044 32160
rect 44060 32096 44124 32160
rect 44140 32096 44204 32160
rect 44220 32096 44284 32160
rect 49740 32156 49804 32160
rect 49820 32156 49884 32160
rect 49740 32100 49754 32156
rect 49754 32100 49804 32156
rect 49820 32100 49834 32156
rect 49834 32100 49884 32156
rect 49740 32096 49804 32100
rect 49820 32096 49884 32100
rect 49900 32096 49964 32160
rect 49980 32096 50044 32160
rect 50060 32096 50124 32160
rect 50140 32096 50204 32160
rect 50220 32096 50284 32160
rect 55740 32096 55804 32160
rect 55820 32096 55884 32160
rect 55900 32096 55964 32160
rect 55980 32096 56044 32160
rect 56060 32096 56124 32160
rect 56140 32096 56204 32160
rect 56220 32096 56284 32160
rect 61740 32096 61804 32160
rect 61820 32096 61884 32160
rect 61900 32096 61964 32160
rect 61980 32096 62044 32160
rect 62060 32096 62124 32160
rect 62140 32096 62204 32160
rect 62220 32096 62284 32160
rect 67740 32096 67804 32160
rect 67820 32096 67884 32160
rect 67900 32096 67964 32160
rect 67980 32096 68044 32160
rect 68060 32096 68124 32160
rect 68140 32096 68204 32160
rect 68220 32096 68284 32160
rect 73740 32096 73804 32160
rect 73820 32096 73884 32160
rect 73900 32096 73964 32160
rect 73980 32096 74044 32160
rect 74060 32096 74124 32160
rect 74140 32096 74204 32160
rect 74220 32096 74284 32160
rect 1740 32016 1804 32080
rect 1820 32016 1884 32080
rect 1900 32016 1964 32080
rect 1980 32016 2044 32080
rect 2060 32016 2124 32080
rect 2140 32016 2204 32080
rect 2220 32076 2284 32080
rect 2220 32020 2276 32076
rect 2276 32020 2284 32076
rect 2220 32016 2284 32020
rect 7740 32016 7804 32080
rect 7820 32016 7884 32080
rect 7900 32016 7964 32080
rect 7980 32016 8044 32080
rect 8060 32016 8124 32080
rect 8140 32016 8204 32080
rect 8220 32016 8284 32080
rect 13740 32016 13804 32080
rect 13820 32016 13884 32080
rect 13900 32016 13964 32080
rect 13980 32016 14044 32080
rect 14060 32016 14124 32080
rect 14140 32076 14204 32080
rect 14140 32020 14155 32076
rect 14155 32020 14204 32076
rect 14140 32016 14204 32020
rect 14220 32016 14284 32080
rect 19740 32016 19804 32080
rect 19820 32016 19884 32080
rect 19900 32076 19964 32080
rect 19980 32076 20044 32080
rect 19900 32020 19935 32076
rect 19935 32020 19964 32076
rect 19980 32020 19991 32076
rect 19991 32020 20044 32076
rect 19900 32016 19964 32020
rect 19980 32016 20044 32020
rect 20060 32016 20124 32080
rect 20140 32016 20204 32080
rect 20220 32016 20284 32080
rect 25740 32076 25804 32080
rect 25740 32020 25771 32076
rect 25771 32020 25804 32076
rect 25740 32016 25804 32020
rect 25820 32016 25884 32080
rect 25900 32016 25964 32080
rect 25980 32016 26044 32080
rect 26060 32016 26124 32080
rect 26140 32016 26204 32080
rect 26220 32016 26284 32080
rect 31740 32016 31804 32080
rect 31820 32016 31884 32080
rect 31900 32016 31964 32080
rect 31980 32016 32044 32080
rect 32060 32016 32124 32080
rect 32140 32016 32204 32080
rect 32220 32016 32284 32080
rect 37740 32016 37804 32080
rect 37820 32016 37884 32080
rect 37900 32016 37964 32080
rect 37980 32016 38044 32080
rect 38060 32016 38124 32080
rect 38140 32016 38204 32080
rect 38220 32016 38284 32080
rect 43740 32016 43804 32080
rect 43820 32016 43884 32080
rect 43900 32016 43964 32080
rect 43980 32016 44044 32080
rect 44060 32016 44124 32080
rect 44140 32016 44204 32080
rect 44220 32016 44284 32080
rect 49740 32076 49804 32080
rect 49820 32076 49884 32080
rect 49740 32020 49754 32076
rect 49754 32020 49804 32076
rect 49820 32020 49834 32076
rect 49834 32020 49884 32076
rect 49740 32016 49804 32020
rect 49820 32016 49884 32020
rect 49900 32016 49964 32080
rect 49980 32016 50044 32080
rect 50060 32016 50124 32080
rect 50140 32016 50204 32080
rect 50220 32016 50284 32080
rect 55740 32016 55804 32080
rect 55820 32016 55884 32080
rect 55900 32016 55964 32080
rect 55980 32016 56044 32080
rect 56060 32016 56124 32080
rect 56140 32016 56204 32080
rect 56220 32016 56284 32080
rect 61740 32016 61804 32080
rect 61820 32016 61884 32080
rect 61900 32016 61964 32080
rect 61980 32016 62044 32080
rect 62060 32016 62124 32080
rect 62140 32016 62204 32080
rect 62220 32016 62284 32080
rect 67740 32016 67804 32080
rect 67820 32016 67884 32080
rect 67900 32016 67964 32080
rect 67980 32016 68044 32080
rect 68060 32016 68124 32080
rect 68140 32016 68204 32080
rect 68220 32016 68284 32080
rect 73740 32016 73804 32080
rect 73820 32016 73884 32080
rect 73900 32016 73964 32080
rect 73980 32016 74044 32080
rect 74060 32016 74124 32080
rect 74140 32016 74204 32080
rect 74220 32016 74284 32080
rect 1740 31936 1804 32000
rect 1820 31936 1884 32000
rect 1900 31936 1964 32000
rect 1980 31936 2044 32000
rect 2060 31936 2124 32000
rect 2140 31936 2204 32000
rect 2220 31996 2284 32000
rect 2220 31940 2276 31996
rect 2276 31940 2284 31996
rect 2220 31936 2284 31940
rect 7740 31936 7804 32000
rect 7820 31936 7884 32000
rect 7900 31936 7964 32000
rect 7980 31936 8044 32000
rect 8060 31936 8124 32000
rect 8140 31936 8204 32000
rect 8220 31936 8284 32000
rect 13740 31936 13804 32000
rect 13820 31936 13884 32000
rect 13900 31936 13964 32000
rect 13980 31936 14044 32000
rect 14060 31936 14124 32000
rect 14140 31996 14204 32000
rect 14140 31940 14155 31996
rect 14155 31940 14204 31996
rect 14140 31936 14204 31940
rect 14220 31936 14284 32000
rect 19740 31936 19804 32000
rect 19820 31936 19884 32000
rect 19900 31996 19964 32000
rect 19980 31996 20044 32000
rect 19900 31940 19935 31996
rect 19935 31940 19964 31996
rect 19980 31940 19991 31996
rect 19991 31940 20044 31996
rect 19900 31936 19964 31940
rect 19980 31936 20044 31940
rect 20060 31936 20124 32000
rect 20140 31936 20204 32000
rect 20220 31936 20284 32000
rect 25740 31996 25804 32000
rect 25740 31940 25771 31996
rect 25771 31940 25804 31996
rect 25740 31936 25804 31940
rect 25820 31936 25884 32000
rect 25900 31936 25964 32000
rect 25980 31936 26044 32000
rect 26060 31936 26124 32000
rect 26140 31936 26204 32000
rect 26220 31936 26284 32000
rect 31740 31936 31804 32000
rect 31820 31936 31884 32000
rect 31900 31936 31964 32000
rect 31980 31936 32044 32000
rect 32060 31936 32124 32000
rect 32140 31936 32204 32000
rect 32220 31936 32284 32000
rect 37740 31936 37804 32000
rect 37820 31936 37884 32000
rect 37900 31936 37964 32000
rect 37980 31936 38044 32000
rect 38060 31936 38124 32000
rect 38140 31936 38204 32000
rect 38220 31936 38284 32000
rect 43740 31936 43804 32000
rect 43820 31936 43884 32000
rect 43900 31936 43964 32000
rect 43980 31936 44044 32000
rect 44060 31936 44124 32000
rect 44140 31936 44204 32000
rect 44220 31936 44284 32000
rect 49740 31996 49804 32000
rect 49820 31996 49884 32000
rect 49740 31940 49754 31996
rect 49754 31940 49804 31996
rect 49820 31940 49834 31996
rect 49834 31940 49884 31996
rect 49740 31936 49804 31940
rect 49820 31936 49884 31940
rect 49900 31936 49964 32000
rect 49980 31936 50044 32000
rect 50060 31936 50124 32000
rect 50140 31936 50204 32000
rect 50220 31936 50284 32000
rect 55740 31936 55804 32000
rect 55820 31936 55884 32000
rect 55900 31936 55964 32000
rect 55980 31936 56044 32000
rect 56060 31936 56124 32000
rect 56140 31936 56204 32000
rect 56220 31936 56284 32000
rect 61740 31936 61804 32000
rect 61820 31936 61884 32000
rect 61900 31936 61964 32000
rect 61980 31936 62044 32000
rect 62060 31936 62124 32000
rect 62140 31936 62204 32000
rect 62220 31936 62284 32000
rect 67740 31936 67804 32000
rect 67820 31936 67884 32000
rect 67900 31936 67964 32000
rect 67980 31936 68044 32000
rect 68060 31936 68124 32000
rect 68140 31936 68204 32000
rect 68220 31936 68284 32000
rect 73740 31936 73804 32000
rect 73820 31936 73884 32000
rect 73900 31936 73964 32000
rect 73980 31936 74044 32000
rect 74060 31936 74124 32000
rect 74140 31936 74204 32000
rect 74220 31936 74284 32000
rect 4740 24528 4804 24592
rect 4820 24528 4884 24592
rect 4900 24528 4964 24592
rect 4980 24528 5044 24592
rect 5060 24528 5124 24592
rect 5140 24528 5204 24592
rect 5220 24528 5284 24592
rect 10740 24528 10804 24592
rect 10820 24528 10884 24592
rect 10900 24528 10964 24592
rect 10980 24528 11044 24592
rect 11060 24528 11124 24592
rect 11140 24528 11204 24592
rect 11220 24528 11284 24592
rect 16740 24528 16804 24592
rect 16820 24528 16884 24592
rect 16900 24528 16964 24592
rect 16980 24528 17044 24592
rect 17060 24528 17124 24592
rect 17140 24588 17204 24592
rect 17220 24588 17284 24592
rect 17140 24532 17192 24588
rect 17192 24532 17204 24588
rect 17220 24532 17248 24588
rect 17248 24532 17284 24588
rect 17140 24528 17204 24532
rect 17220 24528 17284 24532
rect 22740 24528 22804 24592
rect 22820 24528 22884 24592
rect 22900 24528 22964 24592
rect 22980 24588 23044 24592
rect 22980 24532 23028 24588
rect 23028 24532 23044 24588
rect 22980 24528 23044 24532
rect 23060 24528 23124 24592
rect 23140 24528 23204 24592
rect 23220 24528 23284 24592
rect 28740 24588 28804 24592
rect 28740 24532 28752 24588
rect 28752 24532 28804 24588
rect 28740 24528 28804 24532
rect 28820 24528 28884 24592
rect 28900 24528 28964 24592
rect 28980 24528 29044 24592
rect 29060 24528 29124 24592
rect 29140 24528 29204 24592
rect 29220 24528 29284 24592
rect 34740 24528 34804 24592
rect 34820 24528 34884 24592
rect 34900 24528 34964 24592
rect 34980 24528 35044 24592
rect 35060 24528 35124 24592
rect 35140 24528 35204 24592
rect 35220 24528 35284 24592
rect 40740 24528 40804 24592
rect 40820 24528 40884 24592
rect 40900 24528 40964 24592
rect 40980 24528 41044 24592
rect 41060 24528 41124 24592
rect 41140 24528 41204 24592
rect 41220 24528 41284 24592
rect 46740 24528 46804 24592
rect 46820 24528 46884 24592
rect 46900 24528 46964 24592
rect 46980 24528 47044 24592
rect 47060 24528 47124 24592
rect 47140 24528 47204 24592
rect 47220 24528 47284 24592
rect 52740 24528 52804 24592
rect 52820 24528 52884 24592
rect 52900 24528 52964 24592
rect 52980 24528 53044 24592
rect 53060 24528 53124 24592
rect 53140 24528 53204 24592
rect 53220 24528 53284 24592
rect 58740 24528 58804 24592
rect 58820 24528 58884 24592
rect 58900 24528 58964 24592
rect 58980 24528 59044 24592
rect 59060 24528 59124 24592
rect 59140 24588 59204 24592
rect 59140 24532 59196 24588
rect 59196 24532 59204 24588
rect 59140 24528 59204 24532
rect 59220 24528 59284 24592
rect 64740 24528 64804 24592
rect 64820 24528 64884 24592
rect 64900 24528 64964 24592
rect 64980 24528 65044 24592
rect 65060 24528 65124 24592
rect 65140 24528 65204 24592
rect 65220 24528 65284 24592
rect 70740 24528 70804 24592
rect 70820 24528 70884 24592
rect 70900 24528 70964 24592
rect 70980 24528 71044 24592
rect 71060 24528 71124 24592
rect 71140 24528 71204 24592
rect 71220 24528 71284 24592
rect 4740 24448 4804 24512
rect 4820 24448 4884 24512
rect 4900 24448 4964 24512
rect 4980 24448 5044 24512
rect 5060 24448 5124 24512
rect 5140 24448 5204 24512
rect 5220 24448 5284 24512
rect 10740 24448 10804 24512
rect 10820 24448 10884 24512
rect 10900 24448 10964 24512
rect 10980 24448 11044 24512
rect 11060 24448 11124 24512
rect 11140 24448 11204 24512
rect 11220 24448 11284 24512
rect 16740 24448 16804 24512
rect 16820 24448 16884 24512
rect 16900 24448 16964 24512
rect 16980 24448 17044 24512
rect 17060 24448 17124 24512
rect 17140 24508 17204 24512
rect 17220 24508 17284 24512
rect 17140 24452 17192 24508
rect 17192 24452 17204 24508
rect 17220 24452 17248 24508
rect 17248 24452 17284 24508
rect 17140 24448 17204 24452
rect 17220 24448 17284 24452
rect 22740 24448 22804 24512
rect 22820 24448 22884 24512
rect 22900 24448 22964 24512
rect 22980 24508 23044 24512
rect 22980 24452 23028 24508
rect 23028 24452 23044 24508
rect 22980 24448 23044 24452
rect 23060 24448 23124 24512
rect 23140 24448 23204 24512
rect 23220 24448 23284 24512
rect 28740 24508 28804 24512
rect 28740 24452 28752 24508
rect 28752 24452 28804 24508
rect 28740 24448 28804 24452
rect 28820 24448 28884 24512
rect 28900 24448 28964 24512
rect 28980 24448 29044 24512
rect 29060 24448 29124 24512
rect 29140 24448 29204 24512
rect 29220 24448 29284 24512
rect 34740 24448 34804 24512
rect 34820 24448 34884 24512
rect 34900 24448 34964 24512
rect 34980 24448 35044 24512
rect 35060 24448 35124 24512
rect 35140 24448 35204 24512
rect 35220 24448 35284 24512
rect 40740 24448 40804 24512
rect 40820 24448 40884 24512
rect 40900 24448 40964 24512
rect 40980 24448 41044 24512
rect 41060 24448 41124 24512
rect 41140 24448 41204 24512
rect 41220 24448 41284 24512
rect 46740 24448 46804 24512
rect 46820 24448 46884 24512
rect 46900 24448 46964 24512
rect 46980 24448 47044 24512
rect 47060 24448 47124 24512
rect 47140 24448 47204 24512
rect 47220 24448 47284 24512
rect 52740 24448 52804 24512
rect 52820 24448 52884 24512
rect 52900 24448 52964 24512
rect 52980 24448 53044 24512
rect 53060 24448 53124 24512
rect 53140 24448 53204 24512
rect 53220 24448 53284 24512
rect 58740 24448 58804 24512
rect 58820 24448 58884 24512
rect 58900 24448 58964 24512
rect 58980 24448 59044 24512
rect 59060 24448 59124 24512
rect 59140 24508 59204 24512
rect 59140 24452 59196 24508
rect 59196 24452 59204 24508
rect 59140 24448 59204 24452
rect 59220 24448 59284 24512
rect 64740 24448 64804 24512
rect 64820 24448 64884 24512
rect 64900 24448 64964 24512
rect 64980 24448 65044 24512
rect 65060 24448 65124 24512
rect 65140 24448 65204 24512
rect 65220 24448 65284 24512
rect 70740 24448 70804 24512
rect 70820 24448 70884 24512
rect 70900 24448 70964 24512
rect 70980 24448 71044 24512
rect 71060 24448 71124 24512
rect 71140 24448 71204 24512
rect 71220 24448 71284 24512
rect 4740 24368 4804 24432
rect 4820 24368 4884 24432
rect 4900 24368 4964 24432
rect 4980 24368 5044 24432
rect 5060 24368 5124 24432
rect 5140 24368 5204 24432
rect 5220 24368 5284 24432
rect 10740 24368 10804 24432
rect 10820 24368 10884 24432
rect 10900 24368 10964 24432
rect 10980 24368 11044 24432
rect 11060 24368 11124 24432
rect 11140 24368 11204 24432
rect 11220 24368 11284 24432
rect 16740 24368 16804 24432
rect 16820 24368 16884 24432
rect 16900 24368 16964 24432
rect 16980 24368 17044 24432
rect 17060 24368 17124 24432
rect 17140 24428 17204 24432
rect 17220 24428 17284 24432
rect 17140 24372 17192 24428
rect 17192 24372 17204 24428
rect 17220 24372 17248 24428
rect 17248 24372 17284 24428
rect 17140 24368 17204 24372
rect 17220 24368 17284 24372
rect 22740 24368 22804 24432
rect 22820 24368 22884 24432
rect 22900 24368 22964 24432
rect 22980 24428 23044 24432
rect 22980 24372 23028 24428
rect 23028 24372 23044 24428
rect 22980 24368 23044 24372
rect 23060 24368 23124 24432
rect 23140 24368 23204 24432
rect 23220 24368 23284 24432
rect 28740 24428 28804 24432
rect 28740 24372 28752 24428
rect 28752 24372 28804 24428
rect 28740 24368 28804 24372
rect 28820 24368 28884 24432
rect 28900 24368 28964 24432
rect 28980 24368 29044 24432
rect 29060 24368 29124 24432
rect 29140 24368 29204 24432
rect 29220 24368 29284 24432
rect 34740 24368 34804 24432
rect 34820 24368 34884 24432
rect 34900 24368 34964 24432
rect 34980 24368 35044 24432
rect 35060 24368 35124 24432
rect 35140 24368 35204 24432
rect 35220 24368 35284 24432
rect 40740 24368 40804 24432
rect 40820 24368 40884 24432
rect 40900 24368 40964 24432
rect 40980 24368 41044 24432
rect 41060 24368 41124 24432
rect 41140 24368 41204 24432
rect 41220 24368 41284 24432
rect 46740 24368 46804 24432
rect 46820 24368 46884 24432
rect 46900 24368 46964 24432
rect 46980 24368 47044 24432
rect 47060 24368 47124 24432
rect 47140 24368 47204 24432
rect 47220 24368 47284 24432
rect 52740 24368 52804 24432
rect 52820 24368 52884 24432
rect 52900 24368 52964 24432
rect 52980 24368 53044 24432
rect 53060 24368 53124 24432
rect 53140 24368 53204 24432
rect 53220 24368 53284 24432
rect 58740 24368 58804 24432
rect 58820 24368 58884 24432
rect 58900 24368 58964 24432
rect 58980 24368 59044 24432
rect 59060 24368 59124 24432
rect 59140 24428 59204 24432
rect 59140 24372 59196 24428
rect 59196 24372 59204 24428
rect 59140 24368 59204 24372
rect 59220 24368 59284 24432
rect 64740 24368 64804 24432
rect 64820 24368 64884 24432
rect 64900 24368 64964 24432
rect 64980 24368 65044 24432
rect 65060 24368 65124 24432
rect 65140 24368 65204 24432
rect 65220 24368 65284 24432
rect 70740 24368 70804 24432
rect 70820 24368 70884 24432
rect 70900 24368 70964 24432
rect 70980 24368 71044 24432
rect 71060 24368 71124 24432
rect 71140 24368 71204 24432
rect 71220 24368 71284 24432
rect 4740 24288 4804 24352
rect 4820 24288 4884 24352
rect 4900 24288 4964 24352
rect 4980 24288 5044 24352
rect 5060 24288 5124 24352
rect 5140 24288 5204 24352
rect 5220 24288 5284 24352
rect 10740 24288 10804 24352
rect 10820 24288 10884 24352
rect 10900 24288 10964 24352
rect 10980 24288 11044 24352
rect 11060 24288 11124 24352
rect 11140 24288 11204 24352
rect 11220 24288 11284 24352
rect 16740 24288 16804 24352
rect 16820 24288 16884 24352
rect 16900 24288 16964 24352
rect 16980 24288 17044 24352
rect 17060 24288 17124 24352
rect 17140 24348 17204 24352
rect 17220 24348 17284 24352
rect 17140 24292 17192 24348
rect 17192 24292 17204 24348
rect 17220 24292 17248 24348
rect 17248 24292 17284 24348
rect 17140 24288 17204 24292
rect 17220 24288 17284 24292
rect 22740 24288 22804 24352
rect 22820 24288 22884 24352
rect 22900 24288 22964 24352
rect 22980 24348 23044 24352
rect 22980 24292 23028 24348
rect 23028 24292 23044 24348
rect 22980 24288 23044 24292
rect 23060 24288 23124 24352
rect 23140 24288 23204 24352
rect 23220 24288 23284 24352
rect 28740 24348 28804 24352
rect 28740 24292 28752 24348
rect 28752 24292 28804 24348
rect 28740 24288 28804 24292
rect 28820 24288 28884 24352
rect 28900 24288 28964 24352
rect 28980 24288 29044 24352
rect 29060 24288 29124 24352
rect 29140 24288 29204 24352
rect 29220 24288 29284 24352
rect 34740 24288 34804 24352
rect 34820 24288 34884 24352
rect 34900 24288 34964 24352
rect 34980 24288 35044 24352
rect 35060 24288 35124 24352
rect 35140 24288 35204 24352
rect 35220 24288 35284 24352
rect 40740 24288 40804 24352
rect 40820 24288 40884 24352
rect 40900 24288 40964 24352
rect 40980 24288 41044 24352
rect 41060 24288 41124 24352
rect 41140 24288 41204 24352
rect 41220 24288 41284 24352
rect 46740 24288 46804 24352
rect 46820 24288 46884 24352
rect 46900 24288 46964 24352
rect 46980 24288 47044 24352
rect 47060 24288 47124 24352
rect 47140 24288 47204 24352
rect 47220 24288 47284 24352
rect 52740 24288 52804 24352
rect 52820 24288 52884 24352
rect 52900 24288 52964 24352
rect 52980 24288 53044 24352
rect 53060 24288 53124 24352
rect 53140 24288 53204 24352
rect 53220 24288 53284 24352
rect 58740 24288 58804 24352
rect 58820 24288 58884 24352
rect 58900 24288 58964 24352
rect 58980 24288 59044 24352
rect 59060 24288 59124 24352
rect 59140 24348 59204 24352
rect 59140 24292 59196 24348
rect 59196 24292 59204 24348
rect 59140 24288 59204 24292
rect 59220 24288 59284 24352
rect 64740 24288 64804 24352
rect 64820 24288 64884 24352
rect 64900 24288 64964 24352
rect 64980 24288 65044 24352
rect 65060 24288 65124 24352
rect 65140 24288 65204 24352
rect 65220 24288 65284 24352
rect 70740 24288 70804 24352
rect 70820 24288 70884 24352
rect 70900 24288 70964 24352
rect 70980 24288 71044 24352
rect 71060 24288 71124 24352
rect 71140 24288 71204 24352
rect 71220 24288 71284 24352
rect 67036 23564 67100 23628
rect 67220 23488 67284 23492
rect 67220 23432 67270 23488
rect 67270 23432 67284 23488
rect 67220 23428 67284 23432
rect 66484 22672 66548 22676
rect 66484 22616 66534 22672
rect 66534 22616 66548 22672
rect 66484 22612 66548 22616
rect 66300 22400 66364 22404
rect 66300 22344 66314 22400
rect 66314 22344 66364 22400
rect 66300 22340 66364 22344
rect 1740 22176 1804 22240
rect 1820 22176 1884 22240
rect 1900 22176 1964 22240
rect 1980 22176 2044 22240
rect 2060 22176 2124 22240
rect 2140 22176 2204 22240
rect 2220 22236 2284 22240
rect 2220 22180 2276 22236
rect 2276 22180 2284 22236
rect 2220 22176 2284 22180
rect 7740 22176 7804 22240
rect 7820 22176 7884 22240
rect 7900 22176 7964 22240
rect 7980 22176 8044 22240
rect 8060 22176 8124 22240
rect 8140 22176 8204 22240
rect 8220 22176 8284 22240
rect 13740 22176 13804 22240
rect 13820 22176 13884 22240
rect 13900 22176 13964 22240
rect 13980 22176 14044 22240
rect 14060 22176 14124 22240
rect 14140 22236 14204 22240
rect 14140 22180 14155 22236
rect 14155 22180 14204 22236
rect 14140 22176 14204 22180
rect 14220 22176 14284 22240
rect 19740 22176 19804 22240
rect 19820 22176 19884 22240
rect 19900 22236 19964 22240
rect 19980 22236 20044 22240
rect 19900 22180 19935 22236
rect 19935 22180 19964 22236
rect 19980 22180 19991 22236
rect 19991 22180 20044 22236
rect 19900 22176 19964 22180
rect 19980 22176 20044 22180
rect 20060 22176 20124 22240
rect 20140 22176 20204 22240
rect 20220 22176 20284 22240
rect 25740 22236 25804 22240
rect 25740 22180 25771 22236
rect 25771 22180 25804 22236
rect 25740 22176 25804 22180
rect 25820 22176 25884 22240
rect 25900 22176 25964 22240
rect 25980 22176 26044 22240
rect 26060 22176 26124 22240
rect 26140 22176 26204 22240
rect 26220 22176 26284 22240
rect 31740 22176 31804 22240
rect 31820 22176 31884 22240
rect 31900 22176 31964 22240
rect 31980 22176 32044 22240
rect 32060 22176 32124 22240
rect 32140 22176 32204 22240
rect 32220 22176 32284 22240
rect 37740 22176 37804 22240
rect 37820 22176 37884 22240
rect 37900 22176 37964 22240
rect 37980 22176 38044 22240
rect 38060 22176 38124 22240
rect 38140 22176 38204 22240
rect 38220 22176 38284 22240
rect 43740 22176 43804 22240
rect 43820 22176 43884 22240
rect 43900 22176 43964 22240
rect 43980 22176 44044 22240
rect 44060 22176 44124 22240
rect 44140 22176 44204 22240
rect 44220 22176 44284 22240
rect 49740 22236 49804 22240
rect 49820 22236 49884 22240
rect 49740 22180 49754 22236
rect 49754 22180 49804 22236
rect 49820 22180 49834 22236
rect 49834 22180 49884 22236
rect 49740 22176 49804 22180
rect 49820 22176 49884 22180
rect 49900 22176 49964 22240
rect 49980 22176 50044 22240
rect 50060 22176 50124 22240
rect 50140 22176 50204 22240
rect 50220 22176 50284 22240
rect 55740 22176 55804 22240
rect 55820 22176 55884 22240
rect 55900 22176 55964 22240
rect 55980 22176 56044 22240
rect 56060 22176 56124 22240
rect 56140 22176 56204 22240
rect 56220 22176 56284 22240
rect 61740 22176 61804 22240
rect 61820 22176 61884 22240
rect 61900 22176 61964 22240
rect 61980 22176 62044 22240
rect 62060 22176 62124 22240
rect 62140 22176 62204 22240
rect 62220 22176 62284 22240
rect 67740 22176 67804 22240
rect 67820 22176 67884 22240
rect 67900 22176 67964 22240
rect 67980 22176 68044 22240
rect 68060 22176 68124 22240
rect 68140 22176 68204 22240
rect 68220 22176 68284 22240
rect 73740 22176 73804 22240
rect 73820 22176 73884 22240
rect 73900 22176 73964 22240
rect 73980 22176 74044 22240
rect 74060 22176 74124 22240
rect 74140 22176 74204 22240
rect 74220 22176 74284 22240
rect 1740 22096 1804 22160
rect 1820 22096 1884 22160
rect 1900 22096 1964 22160
rect 1980 22096 2044 22160
rect 2060 22096 2124 22160
rect 2140 22096 2204 22160
rect 2220 22156 2284 22160
rect 2220 22100 2276 22156
rect 2276 22100 2284 22156
rect 2220 22096 2284 22100
rect 7740 22096 7804 22160
rect 7820 22096 7884 22160
rect 7900 22096 7964 22160
rect 7980 22096 8044 22160
rect 8060 22096 8124 22160
rect 8140 22096 8204 22160
rect 8220 22096 8284 22160
rect 13740 22096 13804 22160
rect 13820 22096 13884 22160
rect 13900 22096 13964 22160
rect 13980 22096 14044 22160
rect 14060 22096 14124 22160
rect 14140 22156 14204 22160
rect 14140 22100 14155 22156
rect 14155 22100 14204 22156
rect 14140 22096 14204 22100
rect 14220 22096 14284 22160
rect 19740 22096 19804 22160
rect 19820 22096 19884 22160
rect 19900 22156 19964 22160
rect 19980 22156 20044 22160
rect 19900 22100 19935 22156
rect 19935 22100 19964 22156
rect 19980 22100 19991 22156
rect 19991 22100 20044 22156
rect 19900 22096 19964 22100
rect 19980 22096 20044 22100
rect 20060 22096 20124 22160
rect 20140 22096 20204 22160
rect 20220 22096 20284 22160
rect 25740 22156 25804 22160
rect 25740 22100 25771 22156
rect 25771 22100 25804 22156
rect 25740 22096 25804 22100
rect 25820 22096 25884 22160
rect 25900 22096 25964 22160
rect 25980 22096 26044 22160
rect 26060 22096 26124 22160
rect 26140 22096 26204 22160
rect 26220 22096 26284 22160
rect 31740 22096 31804 22160
rect 31820 22096 31884 22160
rect 31900 22096 31964 22160
rect 31980 22096 32044 22160
rect 32060 22096 32124 22160
rect 32140 22096 32204 22160
rect 32220 22096 32284 22160
rect 37740 22096 37804 22160
rect 37820 22096 37884 22160
rect 37900 22096 37964 22160
rect 37980 22096 38044 22160
rect 38060 22096 38124 22160
rect 38140 22096 38204 22160
rect 38220 22096 38284 22160
rect 43740 22096 43804 22160
rect 43820 22096 43884 22160
rect 43900 22096 43964 22160
rect 43980 22096 44044 22160
rect 44060 22096 44124 22160
rect 44140 22096 44204 22160
rect 44220 22096 44284 22160
rect 49740 22156 49804 22160
rect 49820 22156 49884 22160
rect 49740 22100 49754 22156
rect 49754 22100 49804 22156
rect 49820 22100 49834 22156
rect 49834 22100 49884 22156
rect 49740 22096 49804 22100
rect 49820 22096 49884 22100
rect 49900 22096 49964 22160
rect 49980 22096 50044 22160
rect 50060 22096 50124 22160
rect 50140 22096 50204 22160
rect 50220 22096 50284 22160
rect 55740 22096 55804 22160
rect 55820 22096 55884 22160
rect 55900 22096 55964 22160
rect 55980 22096 56044 22160
rect 56060 22096 56124 22160
rect 56140 22096 56204 22160
rect 56220 22096 56284 22160
rect 61740 22096 61804 22160
rect 61820 22096 61884 22160
rect 61900 22096 61964 22160
rect 61980 22096 62044 22160
rect 62060 22096 62124 22160
rect 62140 22096 62204 22160
rect 62220 22096 62284 22160
rect 67740 22096 67804 22160
rect 67820 22096 67884 22160
rect 67900 22096 67964 22160
rect 67980 22096 68044 22160
rect 68060 22096 68124 22160
rect 68140 22096 68204 22160
rect 68220 22096 68284 22160
rect 73740 22096 73804 22160
rect 73820 22096 73884 22160
rect 73900 22096 73964 22160
rect 73980 22096 74044 22160
rect 74060 22096 74124 22160
rect 74140 22096 74204 22160
rect 74220 22096 74284 22160
rect 1740 22016 1804 22080
rect 1820 22016 1884 22080
rect 1900 22016 1964 22080
rect 1980 22016 2044 22080
rect 2060 22016 2124 22080
rect 2140 22016 2204 22080
rect 2220 22076 2284 22080
rect 2220 22020 2276 22076
rect 2276 22020 2284 22076
rect 2220 22016 2284 22020
rect 7740 22016 7804 22080
rect 7820 22016 7884 22080
rect 7900 22016 7964 22080
rect 7980 22016 8044 22080
rect 8060 22016 8124 22080
rect 8140 22016 8204 22080
rect 8220 22016 8284 22080
rect 13740 22016 13804 22080
rect 13820 22016 13884 22080
rect 13900 22016 13964 22080
rect 13980 22016 14044 22080
rect 14060 22016 14124 22080
rect 14140 22076 14204 22080
rect 14140 22020 14155 22076
rect 14155 22020 14204 22076
rect 14140 22016 14204 22020
rect 14220 22016 14284 22080
rect 19740 22016 19804 22080
rect 19820 22016 19884 22080
rect 19900 22076 19964 22080
rect 19980 22076 20044 22080
rect 19900 22020 19935 22076
rect 19935 22020 19964 22076
rect 19980 22020 19991 22076
rect 19991 22020 20044 22076
rect 19900 22016 19964 22020
rect 19980 22016 20044 22020
rect 20060 22016 20124 22080
rect 20140 22016 20204 22080
rect 20220 22016 20284 22080
rect 25740 22076 25804 22080
rect 25740 22020 25771 22076
rect 25771 22020 25804 22076
rect 25740 22016 25804 22020
rect 25820 22016 25884 22080
rect 25900 22016 25964 22080
rect 25980 22016 26044 22080
rect 26060 22016 26124 22080
rect 26140 22016 26204 22080
rect 26220 22016 26284 22080
rect 31740 22016 31804 22080
rect 31820 22016 31884 22080
rect 31900 22016 31964 22080
rect 31980 22016 32044 22080
rect 32060 22016 32124 22080
rect 32140 22016 32204 22080
rect 32220 22016 32284 22080
rect 37740 22016 37804 22080
rect 37820 22016 37884 22080
rect 37900 22016 37964 22080
rect 37980 22016 38044 22080
rect 38060 22016 38124 22080
rect 38140 22016 38204 22080
rect 38220 22016 38284 22080
rect 43740 22016 43804 22080
rect 43820 22016 43884 22080
rect 43900 22016 43964 22080
rect 43980 22016 44044 22080
rect 44060 22016 44124 22080
rect 44140 22016 44204 22080
rect 44220 22016 44284 22080
rect 49740 22076 49804 22080
rect 49820 22076 49884 22080
rect 49740 22020 49754 22076
rect 49754 22020 49804 22076
rect 49820 22020 49834 22076
rect 49834 22020 49884 22076
rect 49740 22016 49804 22020
rect 49820 22016 49884 22020
rect 49900 22016 49964 22080
rect 49980 22016 50044 22080
rect 50060 22016 50124 22080
rect 50140 22016 50204 22080
rect 50220 22016 50284 22080
rect 55740 22016 55804 22080
rect 55820 22016 55884 22080
rect 55900 22016 55964 22080
rect 55980 22016 56044 22080
rect 56060 22016 56124 22080
rect 56140 22016 56204 22080
rect 56220 22016 56284 22080
rect 61740 22016 61804 22080
rect 61820 22016 61884 22080
rect 61900 22016 61964 22080
rect 61980 22016 62044 22080
rect 62060 22016 62124 22080
rect 62140 22016 62204 22080
rect 62220 22016 62284 22080
rect 67740 22016 67804 22080
rect 67820 22016 67884 22080
rect 67900 22016 67964 22080
rect 67980 22016 68044 22080
rect 68060 22016 68124 22080
rect 68140 22016 68204 22080
rect 68220 22016 68284 22080
rect 73740 22016 73804 22080
rect 73820 22016 73884 22080
rect 73900 22016 73964 22080
rect 73980 22016 74044 22080
rect 74060 22016 74124 22080
rect 74140 22016 74204 22080
rect 74220 22016 74284 22080
rect 1740 21936 1804 22000
rect 1820 21936 1884 22000
rect 1900 21936 1964 22000
rect 1980 21936 2044 22000
rect 2060 21936 2124 22000
rect 2140 21936 2204 22000
rect 2220 21996 2284 22000
rect 2220 21940 2276 21996
rect 2276 21940 2284 21996
rect 2220 21936 2284 21940
rect 7740 21936 7804 22000
rect 7820 21936 7884 22000
rect 7900 21936 7964 22000
rect 7980 21936 8044 22000
rect 8060 21936 8124 22000
rect 8140 21936 8204 22000
rect 8220 21936 8284 22000
rect 13740 21936 13804 22000
rect 13820 21936 13884 22000
rect 13900 21936 13964 22000
rect 13980 21936 14044 22000
rect 14060 21936 14124 22000
rect 14140 21996 14204 22000
rect 14140 21940 14155 21996
rect 14155 21940 14204 21996
rect 14140 21936 14204 21940
rect 14220 21936 14284 22000
rect 19740 21936 19804 22000
rect 19820 21936 19884 22000
rect 19900 21996 19964 22000
rect 19980 21996 20044 22000
rect 19900 21940 19935 21996
rect 19935 21940 19964 21996
rect 19980 21940 19991 21996
rect 19991 21940 20044 21996
rect 19900 21936 19964 21940
rect 19980 21936 20044 21940
rect 20060 21936 20124 22000
rect 20140 21936 20204 22000
rect 20220 21936 20284 22000
rect 25740 21996 25804 22000
rect 25740 21940 25771 21996
rect 25771 21940 25804 21996
rect 25740 21936 25804 21940
rect 25820 21936 25884 22000
rect 25900 21936 25964 22000
rect 25980 21936 26044 22000
rect 26060 21936 26124 22000
rect 26140 21936 26204 22000
rect 26220 21936 26284 22000
rect 31740 21936 31804 22000
rect 31820 21936 31884 22000
rect 31900 21936 31964 22000
rect 31980 21936 32044 22000
rect 32060 21936 32124 22000
rect 32140 21936 32204 22000
rect 32220 21936 32284 22000
rect 37740 21936 37804 22000
rect 37820 21936 37884 22000
rect 37900 21936 37964 22000
rect 37980 21936 38044 22000
rect 38060 21936 38124 22000
rect 38140 21936 38204 22000
rect 38220 21936 38284 22000
rect 43740 21936 43804 22000
rect 43820 21936 43884 22000
rect 43900 21936 43964 22000
rect 43980 21936 44044 22000
rect 44060 21936 44124 22000
rect 44140 21936 44204 22000
rect 44220 21936 44284 22000
rect 49740 21996 49804 22000
rect 49820 21996 49884 22000
rect 49740 21940 49754 21996
rect 49754 21940 49804 21996
rect 49820 21940 49834 21996
rect 49834 21940 49884 21996
rect 49740 21936 49804 21940
rect 49820 21936 49884 21940
rect 49900 21936 49964 22000
rect 49980 21936 50044 22000
rect 50060 21936 50124 22000
rect 50140 21936 50204 22000
rect 50220 21936 50284 22000
rect 55740 21936 55804 22000
rect 55820 21936 55884 22000
rect 55900 21936 55964 22000
rect 55980 21936 56044 22000
rect 56060 21936 56124 22000
rect 56140 21936 56204 22000
rect 56220 21936 56284 22000
rect 61740 21936 61804 22000
rect 61820 21936 61884 22000
rect 61900 21936 61964 22000
rect 61980 21936 62044 22000
rect 62060 21936 62124 22000
rect 62140 21936 62204 22000
rect 62220 21936 62284 22000
rect 67740 21936 67804 22000
rect 67820 21936 67884 22000
rect 67900 21936 67964 22000
rect 67980 21936 68044 22000
rect 68060 21936 68124 22000
rect 68140 21936 68204 22000
rect 68220 21936 68284 22000
rect 73740 21936 73804 22000
rect 73820 21936 73884 22000
rect 73900 21936 73964 22000
rect 73980 21936 74044 22000
rect 74060 21936 74124 22000
rect 74140 21936 74204 22000
rect 74220 21936 74284 22000
rect 64460 18124 64524 18188
rect 63172 15812 63236 15876
rect 4740 14528 4804 14592
rect 4820 14528 4884 14592
rect 4900 14528 4964 14592
rect 4980 14528 5044 14592
rect 5060 14528 5124 14592
rect 5140 14528 5204 14592
rect 5220 14528 5284 14592
rect 10740 14528 10804 14592
rect 10820 14528 10884 14592
rect 10900 14528 10964 14592
rect 10980 14528 11044 14592
rect 11060 14528 11124 14592
rect 11140 14528 11204 14592
rect 11220 14528 11284 14592
rect 16740 14528 16804 14592
rect 16820 14528 16884 14592
rect 16900 14528 16964 14592
rect 16980 14528 17044 14592
rect 17060 14528 17124 14592
rect 17140 14588 17204 14592
rect 17220 14588 17284 14592
rect 17140 14532 17192 14588
rect 17192 14532 17204 14588
rect 17220 14532 17248 14588
rect 17248 14532 17284 14588
rect 17140 14528 17204 14532
rect 17220 14528 17284 14532
rect 22740 14528 22804 14592
rect 22820 14528 22884 14592
rect 22900 14528 22964 14592
rect 22980 14588 23044 14592
rect 22980 14532 23028 14588
rect 23028 14532 23044 14588
rect 22980 14528 23044 14532
rect 23060 14528 23124 14592
rect 23140 14528 23204 14592
rect 23220 14528 23284 14592
rect 28740 14588 28804 14592
rect 28740 14532 28752 14588
rect 28752 14532 28804 14588
rect 28740 14528 28804 14532
rect 28820 14528 28884 14592
rect 28900 14528 28964 14592
rect 28980 14528 29044 14592
rect 29060 14528 29124 14592
rect 29140 14528 29204 14592
rect 29220 14528 29284 14592
rect 34740 14528 34804 14592
rect 34820 14528 34884 14592
rect 34900 14528 34964 14592
rect 34980 14528 35044 14592
rect 35060 14528 35124 14592
rect 35140 14528 35204 14592
rect 35220 14528 35284 14592
rect 40740 14528 40804 14592
rect 40820 14528 40884 14592
rect 40900 14528 40964 14592
rect 40980 14528 41044 14592
rect 41060 14528 41124 14592
rect 41140 14528 41204 14592
rect 41220 14528 41284 14592
rect 46740 14528 46804 14592
rect 46820 14528 46884 14592
rect 46900 14528 46964 14592
rect 46980 14528 47044 14592
rect 47060 14528 47124 14592
rect 47140 14528 47204 14592
rect 47220 14528 47284 14592
rect 52740 14528 52804 14592
rect 52820 14528 52884 14592
rect 52900 14528 52964 14592
rect 52980 14528 53044 14592
rect 53060 14528 53124 14592
rect 53140 14528 53204 14592
rect 53220 14528 53284 14592
rect 58740 14528 58804 14592
rect 58820 14528 58884 14592
rect 58900 14528 58964 14592
rect 58980 14528 59044 14592
rect 59060 14528 59124 14592
rect 59140 14588 59204 14592
rect 59140 14532 59196 14588
rect 59196 14532 59204 14588
rect 59140 14528 59204 14532
rect 59220 14528 59284 14592
rect 64740 14528 64804 14592
rect 64820 14528 64884 14592
rect 64900 14528 64964 14592
rect 64980 14528 65044 14592
rect 65060 14528 65124 14592
rect 65140 14528 65204 14592
rect 65220 14528 65284 14592
rect 70740 14528 70804 14592
rect 70820 14528 70884 14592
rect 70900 14528 70964 14592
rect 70980 14528 71044 14592
rect 71060 14528 71124 14592
rect 71140 14528 71204 14592
rect 71220 14528 71284 14592
rect 4740 14448 4804 14512
rect 4820 14448 4884 14512
rect 4900 14448 4964 14512
rect 4980 14448 5044 14512
rect 5060 14448 5124 14512
rect 5140 14448 5204 14512
rect 5220 14448 5284 14512
rect 10740 14448 10804 14512
rect 10820 14448 10884 14512
rect 10900 14448 10964 14512
rect 10980 14448 11044 14512
rect 11060 14448 11124 14512
rect 11140 14448 11204 14512
rect 11220 14448 11284 14512
rect 16740 14448 16804 14512
rect 16820 14448 16884 14512
rect 16900 14448 16964 14512
rect 16980 14448 17044 14512
rect 17060 14448 17124 14512
rect 17140 14508 17204 14512
rect 17220 14508 17284 14512
rect 17140 14452 17192 14508
rect 17192 14452 17204 14508
rect 17220 14452 17248 14508
rect 17248 14452 17284 14508
rect 17140 14448 17204 14452
rect 17220 14448 17284 14452
rect 22740 14448 22804 14512
rect 22820 14448 22884 14512
rect 22900 14448 22964 14512
rect 22980 14508 23044 14512
rect 22980 14452 23028 14508
rect 23028 14452 23044 14508
rect 22980 14448 23044 14452
rect 23060 14448 23124 14512
rect 23140 14448 23204 14512
rect 23220 14448 23284 14512
rect 28740 14508 28804 14512
rect 28740 14452 28752 14508
rect 28752 14452 28804 14508
rect 28740 14448 28804 14452
rect 28820 14448 28884 14512
rect 28900 14448 28964 14512
rect 28980 14448 29044 14512
rect 29060 14448 29124 14512
rect 29140 14448 29204 14512
rect 29220 14448 29284 14512
rect 34740 14448 34804 14512
rect 34820 14448 34884 14512
rect 34900 14448 34964 14512
rect 34980 14448 35044 14512
rect 35060 14448 35124 14512
rect 35140 14448 35204 14512
rect 35220 14448 35284 14512
rect 40740 14448 40804 14512
rect 40820 14448 40884 14512
rect 40900 14448 40964 14512
rect 40980 14448 41044 14512
rect 41060 14448 41124 14512
rect 41140 14448 41204 14512
rect 41220 14448 41284 14512
rect 46740 14448 46804 14512
rect 46820 14448 46884 14512
rect 46900 14448 46964 14512
rect 46980 14448 47044 14512
rect 47060 14448 47124 14512
rect 47140 14448 47204 14512
rect 47220 14448 47284 14512
rect 52740 14448 52804 14512
rect 52820 14448 52884 14512
rect 52900 14448 52964 14512
rect 52980 14448 53044 14512
rect 53060 14448 53124 14512
rect 53140 14448 53204 14512
rect 53220 14448 53284 14512
rect 58740 14448 58804 14512
rect 58820 14448 58884 14512
rect 58900 14448 58964 14512
rect 58980 14448 59044 14512
rect 59060 14448 59124 14512
rect 59140 14508 59204 14512
rect 59140 14452 59196 14508
rect 59196 14452 59204 14508
rect 59140 14448 59204 14452
rect 59220 14448 59284 14512
rect 64740 14448 64804 14512
rect 64820 14448 64884 14512
rect 64900 14448 64964 14512
rect 64980 14448 65044 14512
rect 65060 14448 65124 14512
rect 65140 14448 65204 14512
rect 65220 14448 65284 14512
rect 70740 14448 70804 14512
rect 70820 14448 70884 14512
rect 70900 14448 70964 14512
rect 70980 14448 71044 14512
rect 71060 14448 71124 14512
rect 71140 14448 71204 14512
rect 71220 14448 71284 14512
rect 4740 14368 4804 14432
rect 4820 14368 4884 14432
rect 4900 14368 4964 14432
rect 4980 14368 5044 14432
rect 5060 14368 5124 14432
rect 5140 14368 5204 14432
rect 5220 14368 5284 14432
rect 10740 14368 10804 14432
rect 10820 14368 10884 14432
rect 10900 14368 10964 14432
rect 10980 14368 11044 14432
rect 11060 14368 11124 14432
rect 11140 14368 11204 14432
rect 11220 14368 11284 14432
rect 16740 14368 16804 14432
rect 16820 14368 16884 14432
rect 16900 14368 16964 14432
rect 16980 14368 17044 14432
rect 17060 14368 17124 14432
rect 17140 14428 17204 14432
rect 17220 14428 17284 14432
rect 17140 14372 17192 14428
rect 17192 14372 17204 14428
rect 17220 14372 17248 14428
rect 17248 14372 17284 14428
rect 17140 14368 17204 14372
rect 17220 14368 17284 14372
rect 22740 14368 22804 14432
rect 22820 14368 22884 14432
rect 22900 14368 22964 14432
rect 22980 14428 23044 14432
rect 22980 14372 23028 14428
rect 23028 14372 23044 14428
rect 22980 14368 23044 14372
rect 23060 14368 23124 14432
rect 23140 14368 23204 14432
rect 23220 14368 23284 14432
rect 28740 14428 28804 14432
rect 28740 14372 28752 14428
rect 28752 14372 28804 14428
rect 28740 14368 28804 14372
rect 28820 14368 28884 14432
rect 28900 14368 28964 14432
rect 28980 14368 29044 14432
rect 29060 14368 29124 14432
rect 29140 14368 29204 14432
rect 29220 14368 29284 14432
rect 34740 14368 34804 14432
rect 34820 14368 34884 14432
rect 34900 14368 34964 14432
rect 34980 14368 35044 14432
rect 35060 14368 35124 14432
rect 35140 14368 35204 14432
rect 35220 14368 35284 14432
rect 40740 14368 40804 14432
rect 40820 14368 40884 14432
rect 40900 14368 40964 14432
rect 40980 14368 41044 14432
rect 41060 14368 41124 14432
rect 41140 14368 41204 14432
rect 41220 14368 41284 14432
rect 46740 14368 46804 14432
rect 46820 14368 46884 14432
rect 46900 14368 46964 14432
rect 46980 14368 47044 14432
rect 47060 14368 47124 14432
rect 47140 14368 47204 14432
rect 47220 14368 47284 14432
rect 52740 14368 52804 14432
rect 52820 14368 52884 14432
rect 52900 14368 52964 14432
rect 52980 14368 53044 14432
rect 53060 14368 53124 14432
rect 53140 14368 53204 14432
rect 53220 14368 53284 14432
rect 58740 14368 58804 14432
rect 58820 14368 58884 14432
rect 58900 14368 58964 14432
rect 58980 14368 59044 14432
rect 59060 14368 59124 14432
rect 59140 14428 59204 14432
rect 59140 14372 59196 14428
rect 59196 14372 59204 14428
rect 59140 14368 59204 14372
rect 59220 14368 59284 14432
rect 64740 14368 64804 14432
rect 64820 14368 64884 14432
rect 64900 14368 64964 14432
rect 64980 14368 65044 14432
rect 65060 14368 65124 14432
rect 65140 14368 65204 14432
rect 65220 14368 65284 14432
rect 70740 14368 70804 14432
rect 70820 14368 70884 14432
rect 70900 14368 70964 14432
rect 70980 14368 71044 14432
rect 71060 14368 71124 14432
rect 71140 14368 71204 14432
rect 71220 14368 71284 14432
rect 4740 14288 4804 14352
rect 4820 14288 4884 14352
rect 4900 14288 4964 14352
rect 4980 14288 5044 14352
rect 5060 14288 5124 14352
rect 5140 14288 5204 14352
rect 5220 14288 5284 14352
rect 10740 14288 10804 14352
rect 10820 14288 10884 14352
rect 10900 14288 10964 14352
rect 10980 14288 11044 14352
rect 11060 14288 11124 14352
rect 11140 14288 11204 14352
rect 11220 14288 11284 14352
rect 16740 14288 16804 14352
rect 16820 14288 16884 14352
rect 16900 14288 16964 14352
rect 16980 14288 17044 14352
rect 17060 14288 17124 14352
rect 17140 14348 17204 14352
rect 17220 14348 17284 14352
rect 17140 14292 17192 14348
rect 17192 14292 17204 14348
rect 17220 14292 17248 14348
rect 17248 14292 17284 14348
rect 17140 14288 17204 14292
rect 17220 14288 17284 14292
rect 22740 14288 22804 14352
rect 22820 14288 22884 14352
rect 22900 14288 22964 14352
rect 22980 14348 23044 14352
rect 22980 14292 23028 14348
rect 23028 14292 23044 14348
rect 22980 14288 23044 14292
rect 23060 14288 23124 14352
rect 23140 14288 23204 14352
rect 23220 14288 23284 14352
rect 28740 14348 28804 14352
rect 28740 14292 28752 14348
rect 28752 14292 28804 14348
rect 28740 14288 28804 14292
rect 28820 14288 28884 14352
rect 28900 14288 28964 14352
rect 28980 14288 29044 14352
rect 29060 14288 29124 14352
rect 29140 14288 29204 14352
rect 29220 14288 29284 14352
rect 34740 14288 34804 14352
rect 34820 14288 34884 14352
rect 34900 14288 34964 14352
rect 34980 14288 35044 14352
rect 35060 14288 35124 14352
rect 35140 14288 35204 14352
rect 35220 14288 35284 14352
rect 40740 14288 40804 14352
rect 40820 14288 40884 14352
rect 40900 14288 40964 14352
rect 40980 14288 41044 14352
rect 41060 14288 41124 14352
rect 41140 14288 41204 14352
rect 41220 14288 41284 14352
rect 46740 14288 46804 14352
rect 46820 14288 46884 14352
rect 46900 14288 46964 14352
rect 46980 14288 47044 14352
rect 47060 14288 47124 14352
rect 47140 14288 47204 14352
rect 47220 14288 47284 14352
rect 52740 14288 52804 14352
rect 52820 14288 52884 14352
rect 52900 14288 52964 14352
rect 52980 14288 53044 14352
rect 53060 14288 53124 14352
rect 53140 14288 53204 14352
rect 53220 14288 53284 14352
rect 58740 14288 58804 14352
rect 58820 14288 58884 14352
rect 58900 14288 58964 14352
rect 58980 14288 59044 14352
rect 59060 14288 59124 14352
rect 59140 14348 59204 14352
rect 59140 14292 59196 14348
rect 59196 14292 59204 14348
rect 59140 14288 59204 14292
rect 59220 14288 59284 14352
rect 64740 14288 64804 14352
rect 64820 14288 64884 14352
rect 64900 14288 64964 14352
rect 64980 14288 65044 14352
rect 65060 14288 65124 14352
rect 65140 14288 65204 14352
rect 65220 14288 65284 14352
rect 70740 14288 70804 14352
rect 70820 14288 70884 14352
rect 70900 14288 70964 14352
rect 70980 14288 71044 14352
rect 71060 14288 71124 14352
rect 71140 14288 71204 14352
rect 71220 14288 71284 14352
rect 65932 12684 65996 12748
rect 1740 12176 1804 12240
rect 1820 12176 1884 12240
rect 1900 12176 1964 12240
rect 1980 12176 2044 12240
rect 2060 12176 2124 12240
rect 2140 12176 2204 12240
rect 2220 12236 2284 12240
rect 2220 12180 2276 12236
rect 2276 12180 2284 12236
rect 2220 12176 2284 12180
rect 7740 12176 7804 12240
rect 7820 12176 7884 12240
rect 7900 12176 7964 12240
rect 7980 12176 8044 12240
rect 8060 12176 8124 12240
rect 8140 12176 8204 12240
rect 8220 12176 8284 12240
rect 13740 12176 13804 12240
rect 13820 12176 13884 12240
rect 13900 12176 13964 12240
rect 13980 12176 14044 12240
rect 14060 12176 14124 12240
rect 14140 12236 14204 12240
rect 14140 12180 14155 12236
rect 14155 12180 14204 12236
rect 14140 12176 14204 12180
rect 14220 12176 14284 12240
rect 19740 12176 19804 12240
rect 19820 12176 19884 12240
rect 19900 12236 19964 12240
rect 19980 12236 20044 12240
rect 19900 12180 19935 12236
rect 19935 12180 19964 12236
rect 19980 12180 19991 12236
rect 19991 12180 20044 12236
rect 19900 12176 19964 12180
rect 19980 12176 20044 12180
rect 20060 12176 20124 12240
rect 20140 12176 20204 12240
rect 20220 12176 20284 12240
rect 25740 12236 25804 12240
rect 25740 12180 25771 12236
rect 25771 12180 25804 12236
rect 25740 12176 25804 12180
rect 25820 12176 25884 12240
rect 25900 12176 25964 12240
rect 25980 12176 26044 12240
rect 26060 12176 26124 12240
rect 26140 12176 26204 12240
rect 26220 12176 26284 12240
rect 31740 12176 31804 12240
rect 31820 12176 31884 12240
rect 31900 12176 31964 12240
rect 31980 12176 32044 12240
rect 32060 12176 32124 12240
rect 32140 12176 32204 12240
rect 32220 12176 32284 12240
rect 37740 12176 37804 12240
rect 37820 12176 37884 12240
rect 37900 12176 37964 12240
rect 37980 12176 38044 12240
rect 38060 12176 38124 12240
rect 38140 12176 38204 12240
rect 38220 12176 38284 12240
rect 43740 12176 43804 12240
rect 43820 12176 43884 12240
rect 43900 12176 43964 12240
rect 43980 12176 44044 12240
rect 44060 12176 44124 12240
rect 44140 12176 44204 12240
rect 44220 12176 44284 12240
rect 49740 12236 49804 12240
rect 49820 12236 49884 12240
rect 49740 12180 49754 12236
rect 49754 12180 49804 12236
rect 49820 12180 49834 12236
rect 49834 12180 49884 12236
rect 49740 12176 49804 12180
rect 49820 12176 49884 12180
rect 49900 12176 49964 12240
rect 49980 12176 50044 12240
rect 50060 12176 50124 12240
rect 50140 12176 50204 12240
rect 50220 12176 50284 12240
rect 55740 12176 55804 12240
rect 55820 12176 55884 12240
rect 55900 12176 55964 12240
rect 55980 12176 56044 12240
rect 56060 12176 56124 12240
rect 56140 12176 56204 12240
rect 56220 12176 56284 12240
rect 61740 12176 61804 12240
rect 61820 12176 61884 12240
rect 61900 12176 61964 12240
rect 61980 12176 62044 12240
rect 62060 12176 62124 12240
rect 62140 12176 62204 12240
rect 62220 12176 62284 12240
rect 67740 12176 67804 12240
rect 67820 12176 67884 12240
rect 67900 12176 67964 12240
rect 67980 12176 68044 12240
rect 68060 12176 68124 12240
rect 68140 12176 68204 12240
rect 68220 12176 68284 12240
rect 73740 12176 73804 12240
rect 73820 12176 73884 12240
rect 73900 12176 73964 12240
rect 73980 12176 74044 12240
rect 74060 12176 74124 12240
rect 74140 12176 74204 12240
rect 74220 12176 74284 12240
rect 1740 12096 1804 12160
rect 1820 12096 1884 12160
rect 1900 12096 1964 12160
rect 1980 12096 2044 12160
rect 2060 12096 2124 12160
rect 2140 12096 2204 12160
rect 2220 12156 2284 12160
rect 2220 12100 2276 12156
rect 2276 12100 2284 12156
rect 2220 12096 2284 12100
rect 7740 12096 7804 12160
rect 7820 12096 7884 12160
rect 7900 12096 7964 12160
rect 7980 12096 8044 12160
rect 8060 12096 8124 12160
rect 8140 12096 8204 12160
rect 8220 12096 8284 12160
rect 13740 12096 13804 12160
rect 13820 12096 13884 12160
rect 13900 12096 13964 12160
rect 13980 12096 14044 12160
rect 14060 12096 14124 12160
rect 14140 12156 14204 12160
rect 14140 12100 14155 12156
rect 14155 12100 14204 12156
rect 14140 12096 14204 12100
rect 14220 12096 14284 12160
rect 19740 12096 19804 12160
rect 19820 12096 19884 12160
rect 19900 12156 19964 12160
rect 19980 12156 20044 12160
rect 19900 12100 19935 12156
rect 19935 12100 19964 12156
rect 19980 12100 19991 12156
rect 19991 12100 20044 12156
rect 19900 12096 19964 12100
rect 19980 12096 20044 12100
rect 20060 12096 20124 12160
rect 20140 12096 20204 12160
rect 20220 12096 20284 12160
rect 25740 12156 25804 12160
rect 25740 12100 25771 12156
rect 25771 12100 25804 12156
rect 25740 12096 25804 12100
rect 25820 12096 25884 12160
rect 25900 12096 25964 12160
rect 25980 12096 26044 12160
rect 26060 12096 26124 12160
rect 26140 12096 26204 12160
rect 26220 12096 26284 12160
rect 31740 12096 31804 12160
rect 31820 12096 31884 12160
rect 31900 12096 31964 12160
rect 31980 12096 32044 12160
rect 32060 12096 32124 12160
rect 32140 12096 32204 12160
rect 32220 12096 32284 12160
rect 37740 12096 37804 12160
rect 37820 12096 37884 12160
rect 37900 12096 37964 12160
rect 37980 12096 38044 12160
rect 38060 12096 38124 12160
rect 38140 12096 38204 12160
rect 38220 12096 38284 12160
rect 43740 12096 43804 12160
rect 43820 12096 43884 12160
rect 43900 12096 43964 12160
rect 43980 12096 44044 12160
rect 44060 12096 44124 12160
rect 44140 12096 44204 12160
rect 44220 12096 44284 12160
rect 49740 12156 49804 12160
rect 49820 12156 49884 12160
rect 49740 12100 49754 12156
rect 49754 12100 49804 12156
rect 49820 12100 49834 12156
rect 49834 12100 49884 12156
rect 49740 12096 49804 12100
rect 49820 12096 49884 12100
rect 49900 12096 49964 12160
rect 49980 12096 50044 12160
rect 50060 12096 50124 12160
rect 50140 12096 50204 12160
rect 50220 12096 50284 12160
rect 55740 12096 55804 12160
rect 55820 12096 55884 12160
rect 55900 12096 55964 12160
rect 55980 12096 56044 12160
rect 56060 12096 56124 12160
rect 56140 12096 56204 12160
rect 56220 12096 56284 12160
rect 61740 12096 61804 12160
rect 61820 12096 61884 12160
rect 61900 12096 61964 12160
rect 61980 12096 62044 12160
rect 62060 12096 62124 12160
rect 62140 12096 62204 12160
rect 62220 12096 62284 12160
rect 67740 12096 67804 12160
rect 67820 12096 67884 12160
rect 67900 12096 67964 12160
rect 67980 12096 68044 12160
rect 68060 12096 68124 12160
rect 68140 12096 68204 12160
rect 68220 12096 68284 12160
rect 73740 12096 73804 12160
rect 73820 12096 73884 12160
rect 73900 12096 73964 12160
rect 73980 12096 74044 12160
rect 74060 12096 74124 12160
rect 74140 12096 74204 12160
rect 74220 12096 74284 12160
rect 1740 12016 1804 12080
rect 1820 12016 1884 12080
rect 1900 12016 1964 12080
rect 1980 12016 2044 12080
rect 2060 12016 2124 12080
rect 2140 12016 2204 12080
rect 2220 12076 2284 12080
rect 2220 12020 2276 12076
rect 2276 12020 2284 12076
rect 2220 12016 2284 12020
rect 7740 12016 7804 12080
rect 7820 12016 7884 12080
rect 7900 12016 7964 12080
rect 7980 12016 8044 12080
rect 8060 12016 8124 12080
rect 8140 12016 8204 12080
rect 8220 12016 8284 12080
rect 13740 12016 13804 12080
rect 13820 12016 13884 12080
rect 13900 12016 13964 12080
rect 13980 12016 14044 12080
rect 14060 12016 14124 12080
rect 14140 12076 14204 12080
rect 14140 12020 14155 12076
rect 14155 12020 14204 12076
rect 14140 12016 14204 12020
rect 14220 12016 14284 12080
rect 19740 12016 19804 12080
rect 19820 12016 19884 12080
rect 19900 12076 19964 12080
rect 19980 12076 20044 12080
rect 19900 12020 19935 12076
rect 19935 12020 19964 12076
rect 19980 12020 19991 12076
rect 19991 12020 20044 12076
rect 19900 12016 19964 12020
rect 19980 12016 20044 12020
rect 20060 12016 20124 12080
rect 20140 12016 20204 12080
rect 20220 12016 20284 12080
rect 25740 12076 25804 12080
rect 25740 12020 25771 12076
rect 25771 12020 25804 12076
rect 25740 12016 25804 12020
rect 25820 12016 25884 12080
rect 25900 12016 25964 12080
rect 25980 12016 26044 12080
rect 26060 12016 26124 12080
rect 26140 12016 26204 12080
rect 26220 12016 26284 12080
rect 31740 12016 31804 12080
rect 31820 12016 31884 12080
rect 31900 12016 31964 12080
rect 31980 12016 32044 12080
rect 32060 12016 32124 12080
rect 32140 12016 32204 12080
rect 32220 12016 32284 12080
rect 37740 12016 37804 12080
rect 37820 12016 37884 12080
rect 37900 12016 37964 12080
rect 37980 12016 38044 12080
rect 38060 12016 38124 12080
rect 38140 12016 38204 12080
rect 38220 12016 38284 12080
rect 43740 12016 43804 12080
rect 43820 12016 43884 12080
rect 43900 12016 43964 12080
rect 43980 12016 44044 12080
rect 44060 12016 44124 12080
rect 44140 12016 44204 12080
rect 44220 12016 44284 12080
rect 49740 12076 49804 12080
rect 49820 12076 49884 12080
rect 49740 12020 49754 12076
rect 49754 12020 49804 12076
rect 49820 12020 49834 12076
rect 49834 12020 49884 12076
rect 49740 12016 49804 12020
rect 49820 12016 49884 12020
rect 49900 12016 49964 12080
rect 49980 12016 50044 12080
rect 50060 12016 50124 12080
rect 50140 12016 50204 12080
rect 50220 12016 50284 12080
rect 55740 12016 55804 12080
rect 55820 12016 55884 12080
rect 55900 12016 55964 12080
rect 55980 12016 56044 12080
rect 56060 12016 56124 12080
rect 56140 12016 56204 12080
rect 56220 12016 56284 12080
rect 61740 12016 61804 12080
rect 61820 12016 61884 12080
rect 61900 12016 61964 12080
rect 61980 12016 62044 12080
rect 62060 12016 62124 12080
rect 62140 12016 62204 12080
rect 62220 12016 62284 12080
rect 67740 12016 67804 12080
rect 67820 12016 67884 12080
rect 67900 12016 67964 12080
rect 67980 12016 68044 12080
rect 68060 12016 68124 12080
rect 68140 12016 68204 12080
rect 68220 12016 68284 12080
rect 73740 12016 73804 12080
rect 73820 12016 73884 12080
rect 73900 12016 73964 12080
rect 73980 12016 74044 12080
rect 74060 12016 74124 12080
rect 74140 12016 74204 12080
rect 74220 12016 74284 12080
rect 1740 11936 1804 12000
rect 1820 11936 1884 12000
rect 1900 11936 1964 12000
rect 1980 11936 2044 12000
rect 2060 11936 2124 12000
rect 2140 11936 2204 12000
rect 2220 11996 2284 12000
rect 2220 11940 2276 11996
rect 2276 11940 2284 11996
rect 2220 11936 2284 11940
rect 7740 11936 7804 12000
rect 7820 11936 7884 12000
rect 7900 11936 7964 12000
rect 7980 11936 8044 12000
rect 8060 11936 8124 12000
rect 8140 11936 8204 12000
rect 8220 11936 8284 12000
rect 13740 11936 13804 12000
rect 13820 11936 13884 12000
rect 13900 11936 13964 12000
rect 13980 11936 14044 12000
rect 14060 11936 14124 12000
rect 14140 11996 14204 12000
rect 14140 11940 14155 11996
rect 14155 11940 14204 11996
rect 14140 11936 14204 11940
rect 14220 11936 14284 12000
rect 19740 11936 19804 12000
rect 19820 11936 19884 12000
rect 19900 11996 19964 12000
rect 19980 11996 20044 12000
rect 19900 11940 19935 11996
rect 19935 11940 19964 11996
rect 19980 11940 19991 11996
rect 19991 11940 20044 11996
rect 19900 11936 19964 11940
rect 19980 11936 20044 11940
rect 20060 11936 20124 12000
rect 20140 11936 20204 12000
rect 20220 11936 20284 12000
rect 25740 11996 25804 12000
rect 25740 11940 25771 11996
rect 25771 11940 25804 11996
rect 25740 11936 25804 11940
rect 25820 11936 25884 12000
rect 25900 11936 25964 12000
rect 25980 11936 26044 12000
rect 26060 11936 26124 12000
rect 26140 11936 26204 12000
rect 26220 11936 26284 12000
rect 31740 11936 31804 12000
rect 31820 11936 31884 12000
rect 31900 11936 31964 12000
rect 31980 11936 32044 12000
rect 32060 11936 32124 12000
rect 32140 11936 32204 12000
rect 32220 11936 32284 12000
rect 37740 11936 37804 12000
rect 37820 11936 37884 12000
rect 37900 11936 37964 12000
rect 37980 11936 38044 12000
rect 38060 11936 38124 12000
rect 38140 11936 38204 12000
rect 38220 11936 38284 12000
rect 43740 11936 43804 12000
rect 43820 11936 43884 12000
rect 43900 11936 43964 12000
rect 43980 11936 44044 12000
rect 44060 11936 44124 12000
rect 44140 11936 44204 12000
rect 44220 11936 44284 12000
rect 49740 11996 49804 12000
rect 49820 11996 49884 12000
rect 49740 11940 49754 11996
rect 49754 11940 49804 11996
rect 49820 11940 49834 11996
rect 49834 11940 49884 11996
rect 49740 11936 49804 11940
rect 49820 11936 49884 11940
rect 49900 11936 49964 12000
rect 49980 11936 50044 12000
rect 50060 11936 50124 12000
rect 50140 11936 50204 12000
rect 50220 11936 50284 12000
rect 55740 11936 55804 12000
rect 55820 11936 55884 12000
rect 55900 11936 55964 12000
rect 55980 11936 56044 12000
rect 56060 11936 56124 12000
rect 56140 11936 56204 12000
rect 56220 11936 56284 12000
rect 61740 11936 61804 12000
rect 61820 11936 61884 12000
rect 61900 11936 61964 12000
rect 61980 11936 62044 12000
rect 62060 11936 62124 12000
rect 62140 11936 62204 12000
rect 62220 11936 62284 12000
rect 67740 11936 67804 12000
rect 67820 11936 67884 12000
rect 67900 11936 67964 12000
rect 67980 11936 68044 12000
rect 68060 11936 68124 12000
rect 68140 11936 68204 12000
rect 68220 11936 68284 12000
rect 73740 11936 73804 12000
rect 73820 11936 73884 12000
rect 73900 11936 73964 12000
rect 73980 11936 74044 12000
rect 74060 11936 74124 12000
rect 74140 11936 74204 12000
rect 74220 11936 74284 12000
rect 64460 11732 64524 11796
rect 65932 11732 65996 11796
rect 63356 11460 63420 11524
rect 62988 10508 63052 10572
rect 63356 9964 63420 10028
rect 63172 9828 63236 9892
rect 65748 7788 65812 7852
rect 63540 7516 63604 7580
rect 66116 7380 66180 7444
rect 67036 7244 67100 7308
rect 62988 7108 63052 7172
rect 66300 6972 66364 7036
rect 63908 6700 63972 6764
rect 64276 6564 64340 6628
rect 63724 5884 63788 5948
rect 63356 5476 63420 5540
rect 33916 4856 33980 4860
rect 33916 4800 33966 4856
rect 33966 4800 33980 4856
rect 33916 4796 33980 4800
rect 4740 4528 4804 4592
rect 4820 4528 4884 4592
rect 4900 4528 4964 4592
rect 4980 4528 5044 4592
rect 5060 4528 5124 4592
rect 5140 4528 5204 4592
rect 5220 4528 5284 4592
rect 10740 4528 10804 4592
rect 10820 4528 10884 4592
rect 10900 4528 10964 4592
rect 10980 4528 11044 4592
rect 11060 4528 11124 4592
rect 11140 4528 11204 4592
rect 11220 4528 11284 4592
rect 16740 4528 16804 4592
rect 16820 4528 16884 4592
rect 16900 4528 16964 4592
rect 16980 4528 17044 4592
rect 17060 4528 17124 4592
rect 17140 4528 17204 4592
rect 17220 4528 17284 4592
rect 22740 4528 22804 4592
rect 22820 4528 22884 4592
rect 22900 4528 22964 4592
rect 22980 4528 23044 4592
rect 23060 4528 23124 4592
rect 23140 4528 23204 4592
rect 23220 4528 23284 4592
rect 28740 4528 28804 4592
rect 28820 4528 28884 4592
rect 28900 4528 28964 4592
rect 28980 4528 29044 4592
rect 29060 4528 29124 4592
rect 29140 4528 29204 4592
rect 29220 4528 29284 4592
rect 34740 4528 34804 4592
rect 34820 4528 34884 4592
rect 34900 4528 34964 4592
rect 34980 4528 35044 4592
rect 35060 4528 35124 4592
rect 35140 4528 35204 4592
rect 35220 4528 35284 4592
rect 40740 4528 40804 4592
rect 40820 4528 40884 4592
rect 40900 4528 40964 4592
rect 40980 4528 41044 4592
rect 41060 4528 41124 4592
rect 41140 4528 41204 4592
rect 41220 4528 41284 4592
rect 46740 4528 46804 4592
rect 46820 4528 46884 4592
rect 46900 4528 46964 4592
rect 46980 4528 47044 4592
rect 47060 4528 47124 4592
rect 47140 4528 47204 4592
rect 47220 4528 47284 4592
rect 52740 4528 52804 4592
rect 52820 4528 52884 4592
rect 52900 4528 52964 4592
rect 52980 4528 53044 4592
rect 53060 4528 53124 4592
rect 53140 4528 53204 4592
rect 53220 4528 53284 4592
rect 58740 4528 58804 4592
rect 58820 4528 58884 4592
rect 58900 4528 58964 4592
rect 58980 4528 59044 4592
rect 59060 4528 59124 4592
rect 59140 4528 59204 4592
rect 59220 4528 59284 4592
rect 64740 4528 64804 4592
rect 64820 4528 64884 4592
rect 64900 4528 64964 4592
rect 64980 4528 65044 4592
rect 65060 4528 65124 4592
rect 65140 4528 65204 4592
rect 65220 4528 65284 4592
rect 70740 4528 70804 4592
rect 70820 4528 70884 4592
rect 70900 4528 70964 4592
rect 70980 4528 71044 4592
rect 71060 4528 71124 4592
rect 71140 4528 71204 4592
rect 71220 4528 71284 4592
rect 4740 4448 4804 4512
rect 4820 4448 4884 4512
rect 4900 4448 4964 4512
rect 4980 4448 5044 4512
rect 5060 4448 5124 4512
rect 5140 4448 5204 4512
rect 5220 4448 5284 4512
rect 10740 4448 10804 4512
rect 10820 4448 10884 4512
rect 10900 4448 10964 4512
rect 10980 4448 11044 4512
rect 11060 4448 11124 4512
rect 11140 4448 11204 4512
rect 11220 4448 11284 4512
rect 16740 4448 16804 4512
rect 16820 4448 16884 4512
rect 16900 4448 16964 4512
rect 16980 4448 17044 4512
rect 17060 4448 17124 4512
rect 17140 4448 17204 4512
rect 17220 4448 17284 4512
rect 22740 4448 22804 4512
rect 22820 4448 22884 4512
rect 22900 4448 22964 4512
rect 22980 4448 23044 4512
rect 23060 4448 23124 4512
rect 23140 4448 23204 4512
rect 23220 4448 23284 4512
rect 28740 4448 28804 4512
rect 28820 4448 28884 4512
rect 28900 4448 28964 4512
rect 28980 4448 29044 4512
rect 29060 4448 29124 4512
rect 29140 4448 29204 4512
rect 29220 4448 29284 4512
rect 34740 4448 34804 4512
rect 34820 4448 34884 4512
rect 34900 4448 34964 4512
rect 34980 4448 35044 4512
rect 35060 4448 35124 4512
rect 35140 4448 35204 4512
rect 35220 4448 35284 4512
rect 40740 4448 40804 4512
rect 40820 4448 40884 4512
rect 40900 4448 40964 4512
rect 40980 4448 41044 4512
rect 41060 4448 41124 4512
rect 41140 4448 41204 4512
rect 41220 4448 41284 4512
rect 46740 4448 46804 4512
rect 46820 4448 46884 4512
rect 46900 4448 46964 4512
rect 46980 4448 47044 4512
rect 47060 4448 47124 4512
rect 47140 4448 47204 4512
rect 47220 4448 47284 4512
rect 52740 4448 52804 4512
rect 52820 4448 52884 4512
rect 52900 4448 52964 4512
rect 52980 4448 53044 4512
rect 53060 4448 53124 4512
rect 53140 4448 53204 4512
rect 53220 4448 53284 4512
rect 58740 4448 58804 4512
rect 58820 4448 58884 4512
rect 58900 4448 58964 4512
rect 58980 4448 59044 4512
rect 59060 4448 59124 4512
rect 59140 4448 59204 4512
rect 59220 4448 59284 4512
rect 64740 4448 64804 4512
rect 64820 4448 64884 4512
rect 64900 4448 64964 4512
rect 64980 4448 65044 4512
rect 65060 4448 65124 4512
rect 65140 4448 65204 4512
rect 65220 4448 65284 4512
rect 70740 4448 70804 4512
rect 70820 4448 70884 4512
rect 70900 4448 70964 4512
rect 70980 4448 71044 4512
rect 71060 4448 71124 4512
rect 71140 4448 71204 4512
rect 71220 4448 71284 4512
rect 4740 4368 4804 4432
rect 4820 4368 4884 4432
rect 4900 4368 4964 4432
rect 4980 4368 5044 4432
rect 5060 4368 5124 4432
rect 5140 4368 5204 4432
rect 5220 4368 5284 4432
rect 10740 4368 10804 4432
rect 10820 4368 10884 4432
rect 10900 4368 10964 4432
rect 10980 4368 11044 4432
rect 11060 4368 11124 4432
rect 11140 4368 11204 4432
rect 11220 4368 11284 4432
rect 16740 4368 16804 4432
rect 16820 4368 16884 4432
rect 16900 4368 16964 4432
rect 16980 4368 17044 4432
rect 17060 4368 17124 4432
rect 17140 4368 17204 4432
rect 17220 4368 17284 4432
rect 22740 4368 22804 4432
rect 22820 4368 22884 4432
rect 22900 4368 22964 4432
rect 22980 4368 23044 4432
rect 23060 4368 23124 4432
rect 23140 4368 23204 4432
rect 23220 4368 23284 4432
rect 28740 4368 28804 4432
rect 28820 4368 28884 4432
rect 28900 4368 28964 4432
rect 28980 4368 29044 4432
rect 29060 4368 29124 4432
rect 29140 4368 29204 4432
rect 29220 4368 29284 4432
rect 34740 4368 34804 4432
rect 34820 4368 34884 4432
rect 34900 4368 34964 4432
rect 34980 4368 35044 4432
rect 35060 4368 35124 4432
rect 35140 4368 35204 4432
rect 35220 4368 35284 4432
rect 40740 4368 40804 4432
rect 40820 4368 40884 4432
rect 40900 4368 40964 4432
rect 40980 4368 41044 4432
rect 41060 4368 41124 4432
rect 41140 4368 41204 4432
rect 41220 4368 41284 4432
rect 46740 4368 46804 4432
rect 46820 4368 46884 4432
rect 46900 4368 46964 4432
rect 46980 4368 47044 4432
rect 47060 4368 47124 4432
rect 47140 4368 47204 4432
rect 47220 4368 47284 4432
rect 52740 4368 52804 4432
rect 52820 4368 52884 4432
rect 52900 4368 52964 4432
rect 52980 4368 53044 4432
rect 53060 4368 53124 4432
rect 53140 4368 53204 4432
rect 53220 4368 53284 4432
rect 58740 4368 58804 4432
rect 58820 4368 58884 4432
rect 58900 4368 58964 4432
rect 58980 4368 59044 4432
rect 59060 4368 59124 4432
rect 59140 4368 59204 4432
rect 59220 4368 59284 4432
rect 64740 4368 64804 4432
rect 64820 4368 64884 4432
rect 64900 4368 64964 4432
rect 64980 4368 65044 4432
rect 65060 4368 65124 4432
rect 65140 4368 65204 4432
rect 65220 4368 65284 4432
rect 70740 4368 70804 4432
rect 70820 4368 70884 4432
rect 70900 4368 70964 4432
rect 70980 4368 71044 4432
rect 71060 4368 71124 4432
rect 71140 4368 71204 4432
rect 71220 4368 71284 4432
rect 4740 4288 4804 4352
rect 4820 4288 4884 4352
rect 4900 4288 4964 4352
rect 4980 4288 5044 4352
rect 5060 4288 5124 4352
rect 5140 4288 5204 4352
rect 5220 4288 5284 4352
rect 10740 4288 10804 4352
rect 10820 4288 10884 4352
rect 10900 4288 10964 4352
rect 10980 4288 11044 4352
rect 11060 4288 11124 4352
rect 11140 4288 11204 4352
rect 11220 4288 11284 4352
rect 16740 4288 16804 4352
rect 16820 4288 16884 4352
rect 16900 4288 16964 4352
rect 16980 4288 17044 4352
rect 17060 4288 17124 4352
rect 17140 4288 17204 4352
rect 17220 4288 17284 4352
rect 22740 4288 22804 4352
rect 22820 4288 22884 4352
rect 22900 4288 22964 4352
rect 22980 4288 23044 4352
rect 23060 4288 23124 4352
rect 23140 4288 23204 4352
rect 23220 4288 23284 4352
rect 28740 4288 28804 4352
rect 28820 4288 28884 4352
rect 28900 4288 28964 4352
rect 28980 4288 29044 4352
rect 29060 4288 29124 4352
rect 29140 4288 29204 4352
rect 29220 4288 29284 4352
rect 34740 4288 34804 4352
rect 34820 4288 34884 4352
rect 34900 4288 34964 4352
rect 34980 4288 35044 4352
rect 35060 4288 35124 4352
rect 35140 4288 35204 4352
rect 35220 4288 35284 4352
rect 40740 4288 40804 4352
rect 40820 4288 40884 4352
rect 40900 4288 40964 4352
rect 40980 4288 41044 4352
rect 41060 4288 41124 4352
rect 41140 4288 41204 4352
rect 41220 4288 41284 4352
rect 46740 4288 46804 4352
rect 46820 4288 46884 4352
rect 46900 4288 46964 4352
rect 46980 4288 47044 4352
rect 47060 4288 47124 4352
rect 47140 4288 47204 4352
rect 47220 4288 47284 4352
rect 52740 4288 52804 4352
rect 52820 4288 52884 4352
rect 52900 4288 52964 4352
rect 52980 4288 53044 4352
rect 53060 4288 53124 4352
rect 53140 4288 53204 4352
rect 53220 4288 53284 4352
rect 58740 4288 58804 4352
rect 58820 4288 58884 4352
rect 58900 4288 58964 4352
rect 58980 4288 59044 4352
rect 59060 4288 59124 4352
rect 59140 4288 59204 4352
rect 59220 4288 59284 4352
rect 64740 4288 64804 4352
rect 64820 4288 64884 4352
rect 64900 4288 64964 4352
rect 64980 4288 65044 4352
rect 65060 4288 65124 4352
rect 65140 4288 65204 4352
rect 65220 4288 65284 4352
rect 70740 4288 70804 4352
rect 70820 4288 70884 4352
rect 70900 4288 70964 4352
rect 70980 4288 71044 4352
rect 71060 4288 71124 4352
rect 71140 4288 71204 4352
rect 71220 4288 71284 4352
rect 66484 3844 66548 3908
rect 69060 3708 69124 3772
rect 64092 3300 64156 3364
rect 67220 3028 67284 3092
rect 33916 2544 33980 2548
rect 33916 2488 33930 2544
rect 33930 2488 33980 2544
rect 33916 2484 33980 2488
rect 1740 2176 1804 2240
rect 1820 2236 1884 2240
rect 1900 2236 1964 2240
rect 1980 2236 2044 2240
rect 2060 2236 2124 2240
rect 2140 2236 2204 2240
rect 1820 2180 1864 2236
rect 1864 2180 1884 2236
rect 1900 2180 1920 2236
rect 1920 2180 1944 2236
rect 1944 2180 1964 2236
rect 1980 2180 2000 2236
rect 2000 2180 2024 2236
rect 2024 2180 2044 2236
rect 2060 2180 2080 2236
rect 2080 2180 2104 2236
rect 2104 2180 2124 2236
rect 2140 2180 2160 2236
rect 2160 2180 2204 2236
rect 1820 2176 1884 2180
rect 1900 2176 1964 2180
rect 1980 2176 2044 2180
rect 2060 2176 2124 2180
rect 2140 2176 2204 2180
rect 2220 2176 2284 2240
rect 7740 2176 7804 2240
rect 7820 2176 7884 2240
rect 7900 2176 7964 2240
rect 7980 2176 8044 2240
rect 8060 2176 8124 2240
rect 8140 2176 8204 2240
rect 8220 2176 8284 2240
rect 13740 2176 13804 2240
rect 13820 2176 13884 2240
rect 13900 2176 13964 2240
rect 13980 2176 14044 2240
rect 14060 2176 14124 2240
rect 14140 2176 14204 2240
rect 14220 2176 14284 2240
rect 19740 2176 19804 2240
rect 19820 2176 19884 2240
rect 19900 2176 19964 2240
rect 19980 2176 20044 2240
rect 20060 2176 20124 2240
rect 20140 2176 20204 2240
rect 20220 2176 20284 2240
rect 25740 2176 25804 2240
rect 25820 2176 25884 2240
rect 25900 2176 25964 2240
rect 25980 2176 26044 2240
rect 26060 2176 26124 2240
rect 26140 2176 26204 2240
rect 26220 2176 26284 2240
rect 31740 2176 31804 2240
rect 31820 2236 31884 2240
rect 31900 2236 31964 2240
rect 31980 2236 32044 2240
rect 32060 2236 32124 2240
rect 32140 2236 32204 2240
rect 31820 2180 31864 2236
rect 31864 2180 31884 2236
rect 31900 2180 31920 2236
rect 31920 2180 31944 2236
rect 31944 2180 31964 2236
rect 31980 2180 32000 2236
rect 32000 2180 32024 2236
rect 32024 2180 32044 2236
rect 32060 2180 32080 2236
rect 32080 2180 32104 2236
rect 32104 2180 32124 2236
rect 32140 2180 32160 2236
rect 32160 2180 32204 2236
rect 31820 2176 31884 2180
rect 31900 2176 31964 2180
rect 31980 2176 32044 2180
rect 32060 2176 32124 2180
rect 32140 2176 32204 2180
rect 32220 2176 32284 2240
rect 37740 2176 37804 2240
rect 37820 2176 37884 2240
rect 37900 2176 37964 2240
rect 37980 2176 38044 2240
rect 38060 2176 38124 2240
rect 38140 2176 38204 2240
rect 38220 2176 38284 2240
rect 43740 2176 43804 2240
rect 43820 2176 43884 2240
rect 43900 2176 43964 2240
rect 43980 2176 44044 2240
rect 44060 2176 44124 2240
rect 44140 2176 44204 2240
rect 44220 2176 44284 2240
rect 49740 2176 49804 2240
rect 49820 2176 49884 2240
rect 49900 2176 49964 2240
rect 49980 2176 50044 2240
rect 50060 2176 50124 2240
rect 50140 2176 50204 2240
rect 50220 2176 50284 2240
rect 55740 2176 55804 2240
rect 55820 2176 55884 2240
rect 55900 2176 55964 2240
rect 55980 2176 56044 2240
rect 56060 2176 56124 2240
rect 56140 2176 56204 2240
rect 56220 2176 56284 2240
rect 61740 2176 61804 2240
rect 61820 2236 61884 2240
rect 61900 2236 61964 2240
rect 61980 2236 62044 2240
rect 62060 2236 62124 2240
rect 62140 2236 62204 2240
rect 61820 2180 61864 2236
rect 61864 2180 61884 2236
rect 61900 2180 61920 2236
rect 61920 2180 61944 2236
rect 61944 2180 61964 2236
rect 61980 2180 62000 2236
rect 62000 2180 62024 2236
rect 62024 2180 62044 2236
rect 62060 2180 62080 2236
rect 62080 2180 62104 2236
rect 62104 2180 62124 2236
rect 62140 2180 62160 2236
rect 62160 2180 62204 2236
rect 61820 2176 61884 2180
rect 61900 2176 61964 2180
rect 61980 2176 62044 2180
rect 62060 2176 62124 2180
rect 62140 2176 62204 2180
rect 62220 2176 62284 2240
rect 67740 2176 67804 2240
rect 67820 2176 67884 2240
rect 67900 2176 67964 2240
rect 67980 2176 68044 2240
rect 68060 2176 68124 2240
rect 68140 2176 68204 2240
rect 68220 2176 68284 2240
rect 73740 2176 73804 2240
rect 73820 2176 73884 2240
rect 73900 2176 73964 2240
rect 73980 2176 74044 2240
rect 74060 2176 74124 2240
rect 74140 2176 74204 2240
rect 74220 2176 74284 2240
rect 1740 2096 1804 2160
rect 1820 2156 1884 2160
rect 1900 2156 1964 2160
rect 1980 2156 2044 2160
rect 2060 2156 2124 2160
rect 2140 2156 2204 2160
rect 1820 2100 1864 2156
rect 1864 2100 1884 2156
rect 1900 2100 1920 2156
rect 1920 2100 1944 2156
rect 1944 2100 1964 2156
rect 1980 2100 2000 2156
rect 2000 2100 2024 2156
rect 2024 2100 2044 2156
rect 2060 2100 2080 2156
rect 2080 2100 2104 2156
rect 2104 2100 2124 2156
rect 2140 2100 2160 2156
rect 2160 2100 2204 2156
rect 1820 2096 1884 2100
rect 1900 2096 1964 2100
rect 1980 2096 2044 2100
rect 2060 2096 2124 2100
rect 2140 2096 2204 2100
rect 2220 2096 2284 2160
rect 7740 2096 7804 2160
rect 7820 2096 7884 2160
rect 7900 2096 7964 2160
rect 7980 2096 8044 2160
rect 8060 2096 8124 2160
rect 8140 2096 8204 2160
rect 8220 2096 8284 2160
rect 13740 2096 13804 2160
rect 13820 2096 13884 2160
rect 13900 2096 13964 2160
rect 13980 2096 14044 2160
rect 14060 2096 14124 2160
rect 14140 2096 14204 2160
rect 14220 2096 14284 2160
rect 19740 2096 19804 2160
rect 19820 2096 19884 2160
rect 19900 2096 19964 2160
rect 19980 2096 20044 2160
rect 20060 2096 20124 2160
rect 20140 2096 20204 2160
rect 20220 2096 20284 2160
rect 25740 2096 25804 2160
rect 25820 2096 25884 2160
rect 25900 2096 25964 2160
rect 25980 2096 26044 2160
rect 26060 2096 26124 2160
rect 26140 2096 26204 2160
rect 26220 2096 26284 2160
rect 31740 2096 31804 2160
rect 31820 2156 31884 2160
rect 31900 2156 31964 2160
rect 31980 2156 32044 2160
rect 32060 2156 32124 2160
rect 32140 2156 32204 2160
rect 31820 2100 31864 2156
rect 31864 2100 31884 2156
rect 31900 2100 31920 2156
rect 31920 2100 31944 2156
rect 31944 2100 31964 2156
rect 31980 2100 32000 2156
rect 32000 2100 32024 2156
rect 32024 2100 32044 2156
rect 32060 2100 32080 2156
rect 32080 2100 32104 2156
rect 32104 2100 32124 2156
rect 32140 2100 32160 2156
rect 32160 2100 32204 2156
rect 31820 2096 31884 2100
rect 31900 2096 31964 2100
rect 31980 2096 32044 2100
rect 32060 2096 32124 2100
rect 32140 2096 32204 2100
rect 32220 2096 32284 2160
rect 37740 2096 37804 2160
rect 37820 2096 37884 2160
rect 37900 2096 37964 2160
rect 37980 2096 38044 2160
rect 38060 2096 38124 2160
rect 38140 2096 38204 2160
rect 38220 2096 38284 2160
rect 43740 2096 43804 2160
rect 43820 2096 43884 2160
rect 43900 2096 43964 2160
rect 43980 2096 44044 2160
rect 44060 2096 44124 2160
rect 44140 2096 44204 2160
rect 44220 2096 44284 2160
rect 49740 2096 49804 2160
rect 49820 2096 49884 2160
rect 49900 2096 49964 2160
rect 49980 2096 50044 2160
rect 50060 2096 50124 2160
rect 50140 2096 50204 2160
rect 50220 2096 50284 2160
rect 55740 2096 55804 2160
rect 55820 2096 55884 2160
rect 55900 2096 55964 2160
rect 55980 2096 56044 2160
rect 56060 2096 56124 2160
rect 56140 2096 56204 2160
rect 56220 2096 56284 2160
rect 61740 2096 61804 2160
rect 61820 2156 61884 2160
rect 61900 2156 61964 2160
rect 61980 2156 62044 2160
rect 62060 2156 62124 2160
rect 62140 2156 62204 2160
rect 61820 2100 61864 2156
rect 61864 2100 61884 2156
rect 61900 2100 61920 2156
rect 61920 2100 61944 2156
rect 61944 2100 61964 2156
rect 61980 2100 62000 2156
rect 62000 2100 62024 2156
rect 62024 2100 62044 2156
rect 62060 2100 62080 2156
rect 62080 2100 62104 2156
rect 62104 2100 62124 2156
rect 62140 2100 62160 2156
rect 62160 2100 62204 2156
rect 61820 2096 61884 2100
rect 61900 2096 61964 2100
rect 61980 2096 62044 2100
rect 62060 2096 62124 2100
rect 62140 2096 62204 2100
rect 62220 2096 62284 2160
rect 67740 2096 67804 2160
rect 67820 2096 67884 2160
rect 67900 2096 67964 2160
rect 67980 2096 68044 2160
rect 68060 2096 68124 2160
rect 68140 2096 68204 2160
rect 68220 2096 68284 2160
rect 73740 2096 73804 2160
rect 73820 2096 73884 2160
rect 73900 2096 73964 2160
rect 73980 2096 74044 2160
rect 74060 2096 74124 2160
rect 74140 2096 74204 2160
rect 74220 2096 74284 2160
rect 1740 2016 1804 2080
rect 1820 2076 1884 2080
rect 1900 2076 1964 2080
rect 1980 2076 2044 2080
rect 2060 2076 2124 2080
rect 2140 2076 2204 2080
rect 1820 2020 1864 2076
rect 1864 2020 1884 2076
rect 1900 2020 1920 2076
rect 1920 2020 1944 2076
rect 1944 2020 1964 2076
rect 1980 2020 2000 2076
rect 2000 2020 2024 2076
rect 2024 2020 2044 2076
rect 2060 2020 2080 2076
rect 2080 2020 2104 2076
rect 2104 2020 2124 2076
rect 2140 2020 2160 2076
rect 2160 2020 2204 2076
rect 1820 2016 1884 2020
rect 1900 2016 1964 2020
rect 1980 2016 2044 2020
rect 2060 2016 2124 2020
rect 2140 2016 2204 2020
rect 2220 2016 2284 2080
rect 7740 2016 7804 2080
rect 7820 2016 7884 2080
rect 7900 2016 7964 2080
rect 7980 2016 8044 2080
rect 8060 2016 8124 2080
rect 8140 2016 8204 2080
rect 8220 2016 8284 2080
rect 13740 2016 13804 2080
rect 13820 2016 13884 2080
rect 13900 2016 13964 2080
rect 13980 2016 14044 2080
rect 14060 2016 14124 2080
rect 14140 2016 14204 2080
rect 14220 2016 14284 2080
rect 19740 2016 19804 2080
rect 19820 2016 19884 2080
rect 19900 2016 19964 2080
rect 19980 2016 20044 2080
rect 20060 2016 20124 2080
rect 20140 2016 20204 2080
rect 20220 2016 20284 2080
rect 25740 2016 25804 2080
rect 25820 2016 25884 2080
rect 25900 2016 25964 2080
rect 25980 2016 26044 2080
rect 26060 2016 26124 2080
rect 26140 2016 26204 2080
rect 26220 2016 26284 2080
rect 31740 2016 31804 2080
rect 31820 2076 31884 2080
rect 31900 2076 31964 2080
rect 31980 2076 32044 2080
rect 32060 2076 32124 2080
rect 32140 2076 32204 2080
rect 31820 2020 31864 2076
rect 31864 2020 31884 2076
rect 31900 2020 31920 2076
rect 31920 2020 31944 2076
rect 31944 2020 31964 2076
rect 31980 2020 32000 2076
rect 32000 2020 32024 2076
rect 32024 2020 32044 2076
rect 32060 2020 32080 2076
rect 32080 2020 32104 2076
rect 32104 2020 32124 2076
rect 32140 2020 32160 2076
rect 32160 2020 32204 2076
rect 31820 2016 31884 2020
rect 31900 2016 31964 2020
rect 31980 2016 32044 2020
rect 32060 2016 32124 2020
rect 32140 2016 32204 2020
rect 32220 2016 32284 2080
rect 37740 2016 37804 2080
rect 37820 2016 37884 2080
rect 37900 2016 37964 2080
rect 37980 2016 38044 2080
rect 38060 2016 38124 2080
rect 38140 2016 38204 2080
rect 38220 2016 38284 2080
rect 43740 2016 43804 2080
rect 43820 2016 43884 2080
rect 43900 2016 43964 2080
rect 43980 2016 44044 2080
rect 44060 2016 44124 2080
rect 44140 2016 44204 2080
rect 44220 2016 44284 2080
rect 49740 2016 49804 2080
rect 49820 2016 49884 2080
rect 49900 2016 49964 2080
rect 49980 2016 50044 2080
rect 50060 2016 50124 2080
rect 50140 2016 50204 2080
rect 50220 2016 50284 2080
rect 55740 2016 55804 2080
rect 55820 2016 55884 2080
rect 55900 2016 55964 2080
rect 55980 2016 56044 2080
rect 56060 2016 56124 2080
rect 56140 2016 56204 2080
rect 56220 2016 56284 2080
rect 61740 2016 61804 2080
rect 61820 2076 61884 2080
rect 61900 2076 61964 2080
rect 61980 2076 62044 2080
rect 62060 2076 62124 2080
rect 62140 2076 62204 2080
rect 61820 2020 61864 2076
rect 61864 2020 61884 2076
rect 61900 2020 61920 2076
rect 61920 2020 61944 2076
rect 61944 2020 61964 2076
rect 61980 2020 62000 2076
rect 62000 2020 62024 2076
rect 62024 2020 62044 2076
rect 62060 2020 62080 2076
rect 62080 2020 62104 2076
rect 62104 2020 62124 2076
rect 62140 2020 62160 2076
rect 62160 2020 62204 2076
rect 61820 2016 61884 2020
rect 61900 2016 61964 2020
rect 61980 2016 62044 2020
rect 62060 2016 62124 2020
rect 62140 2016 62204 2020
rect 62220 2016 62284 2080
rect 67740 2016 67804 2080
rect 67820 2016 67884 2080
rect 67900 2016 67964 2080
rect 67980 2016 68044 2080
rect 68060 2016 68124 2080
rect 68140 2016 68204 2080
rect 68220 2016 68284 2080
rect 73740 2016 73804 2080
rect 73820 2016 73884 2080
rect 73900 2016 73964 2080
rect 73980 2016 74044 2080
rect 74060 2016 74124 2080
rect 74140 2016 74204 2080
rect 74220 2016 74284 2080
rect 1740 1936 1804 2000
rect 1820 1996 1884 2000
rect 1900 1996 1964 2000
rect 1980 1996 2044 2000
rect 2060 1996 2124 2000
rect 2140 1996 2204 2000
rect 1820 1940 1864 1996
rect 1864 1940 1884 1996
rect 1900 1940 1920 1996
rect 1920 1940 1944 1996
rect 1944 1940 1964 1996
rect 1980 1940 2000 1996
rect 2000 1940 2024 1996
rect 2024 1940 2044 1996
rect 2060 1940 2080 1996
rect 2080 1940 2104 1996
rect 2104 1940 2124 1996
rect 2140 1940 2160 1996
rect 2160 1940 2204 1996
rect 1820 1936 1884 1940
rect 1900 1936 1964 1940
rect 1980 1936 2044 1940
rect 2060 1936 2124 1940
rect 2140 1936 2204 1940
rect 2220 1936 2284 2000
rect 7740 1936 7804 2000
rect 7820 1936 7884 2000
rect 7900 1936 7964 2000
rect 7980 1936 8044 2000
rect 8060 1936 8124 2000
rect 8140 1936 8204 2000
rect 8220 1936 8284 2000
rect 13740 1936 13804 2000
rect 13820 1936 13884 2000
rect 13900 1936 13964 2000
rect 13980 1936 14044 2000
rect 14060 1936 14124 2000
rect 14140 1936 14204 2000
rect 14220 1936 14284 2000
rect 19740 1936 19804 2000
rect 19820 1936 19884 2000
rect 19900 1936 19964 2000
rect 19980 1936 20044 2000
rect 20060 1936 20124 2000
rect 20140 1936 20204 2000
rect 20220 1936 20284 2000
rect 25740 1936 25804 2000
rect 25820 1936 25884 2000
rect 25900 1936 25964 2000
rect 25980 1936 26044 2000
rect 26060 1936 26124 2000
rect 26140 1936 26204 2000
rect 26220 1936 26284 2000
rect 31740 1936 31804 2000
rect 31820 1996 31884 2000
rect 31900 1996 31964 2000
rect 31980 1996 32044 2000
rect 32060 1996 32124 2000
rect 32140 1996 32204 2000
rect 31820 1940 31864 1996
rect 31864 1940 31884 1996
rect 31900 1940 31920 1996
rect 31920 1940 31944 1996
rect 31944 1940 31964 1996
rect 31980 1940 32000 1996
rect 32000 1940 32024 1996
rect 32024 1940 32044 1996
rect 32060 1940 32080 1996
rect 32080 1940 32104 1996
rect 32104 1940 32124 1996
rect 32140 1940 32160 1996
rect 32160 1940 32204 1996
rect 31820 1936 31884 1940
rect 31900 1936 31964 1940
rect 31980 1936 32044 1940
rect 32060 1936 32124 1940
rect 32140 1936 32204 1940
rect 32220 1936 32284 2000
rect 37740 1936 37804 2000
rect 37820 1936 37884 2000
rect 37900 1936 37964 2000
rect 37980 1936 38044 2000
rect 38060 1936 38124 2000
rect 38140 1936 38204 2000
rect 38220 1936 38284 2000
rect 43740 1936 43804 2000
rect 43820 1936 43884 2000
rect 43900 1936 43964 2000
rect 43980 1936 44044 2000
rect 44060 1936 44124 2000
rect 44140 1936 44204 2000
rect 44220 1936 44284 2000
rect 49740 1936 49804 2000
rect 49820 1936 49884 2000
rect 49900 1936 49964 2000
rect 49980 1936 50044 2000
rect 50060 1936 50124 2000
rect 50140 1936 50204 2000
rect 50220 1936 50284 2000
rect 55740 1936 55804 2000
rect 55820 1936 55884 2000
rect 55900 1936 55964 2000
rect 55980 1936 56044 2000
rect 56060 1936 56124 2000
rect 56140 1936 56204 2000
rect 56220 1936 56284 2000
rect 61740 1936 61804 2000
rect 61820 1996 61884 2000
rect 61900 1996 61964 2000
rect 61980 1996 62044 2000
rect 62060 1996 62124 2000
rect 62140 1996 62204 2000
rect 61820 1940 61864 1996
rect 61864 1940 61884 1996
rect 61900 1940 61920 1996
rect 61920 1940 61944 1996
rect 61944 1940 61964 1996
rect 61980 1940 62000 1996
rect 62000 1940 62024 1996
rect 62024 1940 62044 1996
rect 62060 1940 62080 1996
rect 62080 1940 62104 1996
rect 62104 1940 62124 1996
rect 62140 1940 62160 1996
rect 62160 1940 62204 1996
rect 61820 1936 61884 1940
rect 61900 1936 61964 1940
rect 61980 1936 62044 1940
rect 62060 1936 62124 1940
rect 62140 1936 62204 1940
rect 62220 1936 62284 2000
rect 67740 1936 67804 2000
rect 67820 1936 67884 2000
rect 67900 1936 67964 2000
rect 67980 1936 68044 2000
rect 68060 1936 68124 2000
rect 68140 1936 68204 2000
rect 68220 1936 68284 2000
rect 73740 1936 73804 2000
rect 73820 1936 73884 2000
rect 73900 1936 73964 2000
rect 73980 1936 74044 2000
rect 74060 1936 74124 2000
rect 74140 1936 74204 2000
rect 74220 1936 74284 2000
rect 65564 1260 65628 1324
<< metal4 >>
rect 1702 82240 2322 87000
rect 1702 82176 1740 82240
rect 1804 82176 1820 82240
rect 1884 82176 1900 82240
rect 1964 82176 1980 82240
rect 2044 82176 2060 82240
rect 2124 82176 2140 82240
rect 2204 82176 2220 82240
rect 2284 82176 2322 82240
rect 1702 82160 2322 82176
rect 1702 82096 1740 82160
rect 1804 82096 1820 82160
rect 1884 82096 1900 82160
rect 1964 82096 1980 82160
rect 2044 82096 2060 82160
rect 2124 82096 2140 82160
rect 2204 82096 2220 82160
rect 2284 82096 2322 82160
rect 1702 82080 2322 82096
rect 1702 82016 1740 82080
rect 1804 82016 1820 82080
rect 1884 82016 1900 82080
rect 1964 82016 1980 82080
rect 2044 82016 2060 82080
rect 2124 82016 2140 82080
rect 2204 82016 2220 82080
rect 2284 82016 2322 82080
rect 1702 82000 2322 82016
rect 1702 81936 1740 82000
rect 1804 81936 1820 82000
rect 1884 81936 1900 82000
rect 1964 81936 1980 82000
rect 2044 81936 2060 82000
rect 2124 81936 2140 82000
rect 2204 81936 2220 82000
rect 2284 81936 2322 82000
rect 1702 72240 2322 81936
rect 1702 72176 1740 72240
rect 1804 72176 1820 72240
rect 1884 72176 1900 72240
rect 1964 72176 1980 72240
rect 2044 72176 2060 72240
rect 2124 72176 2140 72240
rect 2204 72176 2220 72240
rect 2284 72176 2322 72240
rect 1702 72160 2322 72176
rect 1702 72096 1740 72160
rect 1804 72096 1820 72160
rect 1884 72096 1900 72160
rect 1964 72096 1980 72160
rect 2044 72096 2060 72160
rect 2124 72096 2140 72160
rect 2204 72096 2220 72160
rect 2284 72096 2322 72160
rect 1702 72080 2322 72096
rect 1702 72016 1740 72080
rect 1804 72016 1820 72080
rect 1884 72016 1900 72080
rect 1964 72016 1980 72080
rect 2044 72016 2060 72080
rect 2124 72016 2140 72080
rect 2204 72016 2220 72080
rect 2284 72016 2322 72080
rect 1702 72000 2322 72016
rect 1702 71936 1740 72000
rect 1804 71936 1820 72000
rect 1884 71936 1900 72000
rect 1964 71936 1980 72000
rect 2044 71936 2060 72000
rect 2124 71936 2140 72000
rect 2204 71936 2220 72000
rect 2284 71936 2322 72000
rect 1702 62240 2322 71936
rect 1702 62176 1740 62240
rect 1804 62176 1820 62240
rect 1884 62176 1900 62240
rect 1964 62176 1980 62240
rect 2044 62176 2060 62240
rect 2124 62176 2140 62240
rect 2204 62176 2220 62240
rect 2284 62176 2322 62240
rect 1702 62160 2322 62176
rect 1702 62096 1740 62160
rect 1804 62096 1820 62160
rect 1884 62096 1900 62160
rect 1964 62096 1980 62160
rect 2044 62096 2060 62160
rect 2124 62096 2140 62160
rect 2204 62096 2220 62160
rect 2284 62096 2322 62160
rect 1702 62080 2322 62096
rect 1702 62016 1740 62080
rect 1804 62016 1820 62080
rect 1884 62016 1900 62080
rect 1964 62016 1980 62080
rect 2044 62016 2060 62080
rect 2124 62016 2140 62080
rect 2204 62016 2220 62080
rect 2284 62016 2322 62080
rect 1702 62000 2322 62016
rect 1702 61936 1740 62000
rect 1804 61936 1820 62000
rect 1884 61936 1900 62000
rect 1964 61936 1980 62000
rect 2044 61936 2060 62000
rect 2124 61936 2140 62000
rect 2204 61936 2220 62000
rect 2284 61936 2322 62000
rect 1702 52240 2322 61936
rect 1702 52176 1740 52240
rect 1804 52176 1820 52240
rect 1884 52176 1900 52240
rect 1964 52176 1980 52240
rect 2044 52176 2060 52240
rect 2124 52176 2140 52240
rect 2204 52176 2220 52240
rect 2284 52176 2322 52240
rect 1702 52160 2322 52176
rect 1702 52096 1740 52160
rect 1804 52096 1820 52160
rect 1884 52096 1900 52160
rect 1964 52096 1980 52160
rect 2044 52096 2060 52160
rect 2124 52096 2140 52160
rect 2204 52096 2220 52160
rect 2284 52096 2322 52160
rect 1702 52080 2322 52096
rect 1702 52016 1740 52080
rect 1804 52016 1820 52080
rect 1884 52016 1900 52080
rect 1964 52016 1980 52080
rect 2044 52016 2060 52080
rect 2124 52016 2140 52080
rect 2204 52016 2220 52080
rect 2284 52016 2322 52080
rect 1702 52000 2322 52016
rect 1702 51936 1740 52000
rect 1804 51936 1820 52000
rect 1884 51936 1900 52000
rect 1964 51936 1980 52000
rect 2044 51936 2060 52000
rect 2124 51936 2140 52000
rect 2204 51936 2220 52000
rect 2284 51936 2322 52000
rect 1702 42240 2322 51936
rect 1702 42176 1740 42240
rect 1804 42176 1820 42240
rect 1884 42176 1900 42240
rect 1964 42176 1980 42240
rect 2044 42176 2060 42240
rect 2124 42176 2140 42240
rect 2204 42176 2220 42240
rect 2284 42176 2322 42240
rect 1702 42160 2322 42176
rect 1702 42096 1740 42160
rect 1804 42096 1820 42160
rect 1884 42096 1900 42160
rect 1964 42096 1980 42160
rect 2044 42096 2060 42160
rect 2124 42096 2140 42160
rect 2204 42096 2220 42160
rect 2284 42096 2322 42160
rect 1702 42080 2322 42096
rect 1702 42016 1740 42080
rect 1804 42016 1820 42080
rect 1884 42016 1900 42080
rect 1964 42016 1980 42080
rect 2044 42016 2060 42080
rect 2124 42016 2140 42080
rect 2204 42016 2220 42080
rect 2284 42016 2322 42080
rect 1702 42000 2322 42016
rect 1702 41936 1740 42000
rect 1804 41936 1820 42000
rect 1884 41936 1900 42000
rect 1964 41936 1980 42000
rect 2044 41936 2060 42000
rect 2124 41936 2140 42000
rect 2204 41936 2220 42000
rect 2284 41936 2322 42000
rect 1702 32240 2322 41936
rect 1702 32176 1740 32240
rect 1804 32176 1820 32240
rect 1884 32176 1900 32240
rect 1964 32176 1980 32240
rect 2044 32176 2060 32240
rect 2124 32176 2140 32240
rect 2204 32176 2220 32240
rect 2284 32176 2322 32240
rect 1702 32160 2322 32176
rect 1702 32096 1740 32160
rect 1804 32096 1820 32160
rect 1884 32096 1900 32160
rect 1964 32096 1980 32160
rect 2044 32096 2060 32160
rect 2124 32096 2140 32160
rect 2204 32096 2220 32160
rect 2284 32096 2322 32160
rect 1702 32080 2322 32096
rect 1702 32016 1740 32080
rect 1804 32016 1820 32080
rect 1884 32016 1900 32080
rect 1964 32016 1980 32080
rect 2044 32016 2060 32080
rect 2124 32016 2140 32080
rect 2204 32016 2220 32080
rect 2284 32016 2322 32080
rect 1702 32000 2322 32016
rect 1702 31936 1740 32000
rect 1804 31936 1820 32000
rect 1884 31936 1900 32000
rect 1964 31936 1980 32000
rect 2044 31936 2060 32000
rect 2124 31936 2140 32000
rect 2204 31936 2220 32000
rect 2284 31936 2322 32000
rect 1702 22240 2322 31936
rect 1702 22176 1740 22240
rect 1804 22176 1820 22240
rect 1884 22176 1900 22240
rect 1964 22176 1980 22240
rect 2044 22176 2060 22240
rect 2124 22176 2140 22240
rect 2204 22176 2220 22240
rect 2284 22176 2322 22240
rect 1702 22160 2322 22176
rect 1702 22096 1740 22160
rect 1804 22096 1820 22160
rect 1884 22096 1900 22160
rect 1964 22096 1980 22160
rect 2044 22096 2060 22160
rect 2124 22096 2140 22160
rect 2204 22096 2220 22160
rect 2284 22096 2322 22160
rect 1702 22080 2322 22096
rect 1702 22016 1740 22080
rect 1804 22016 1820 22080
rect 1884 22016 1900 22080
rect 1964 22016 1980 22080
rect 2044 22016 2060 22080
rect 2124 22016 2140 22080
rect 2204 22016 2220 22080
rect 2284 22016 2322 22080
rect 1702 22000 2322 22016
rect 1702 21936 1740 22000
rect 1804 21936 1820 22000
rect 1884 21936 1900 22000
rect 1964 21936 1980 22000
rect 2044 21936 2060 22000
rect 2124 21936 2140 22000
rect 2204 21936 2220 22000
rect 2284 21936 2322 22000
rect 1702 12240 2322 21936
rect 1702 12176 1740 12240
rect 1804 12176 1820 12240
rect 1884 12176 1900 12240
rect 1964 12176 1980 12240
rect 2044 12176 2060 12240
rect 2124 12176 2140 12240
rect 2204 12176 2220 12240
rect 2284 12176 2322 12240
rect 1702 12160 2322 12176
rect 1702 12096 1740 12160
rect 1804 12096 1820 12160
rect 1884 12096 1900 12160
rect 1964 12096 1980 12160
rect 2044 12096 2060 12160
rect 2124 12096 2140 12160
rect 2204 12096 2220 12160
rect 2284 12096 2322 12160
rect 1702 12080 2322 12096
rect 1702 12016 1740 12080
rect 1804 12016 1820 12080
rect 1884 12016 1900 12080
rect 1964 12016 1980 12080
rect 2044 12016 2060 12080
rect 2124 12016 2140 12080
rect 2204 12016 2220 12080
rect 2284 12016 2322 12080
rect 1702 12000 2322 12016
rect 1702 11936 1740 12000
rect 1804 11936 1820 12000
rect 1884 11936 1900 12000
rect 1964 11936 1980 12000
rect 2044 11936 2060 12000
rect 2124 11936 2140 12000
rect 2204 11936 2220 12000
rect 2284 11936 2322 12000
rect 1702 2240 2322 11936
rect 1702 2176 1740 2240
rect 1804 2176 1820 2240
rect 1884 2176 1900 2240
rect 1964 2176 1980 2240
rect 2044 2176 2060 2240
rect 2124 2176 2140 2240
rect 2204 2176 2220 2240
rect 2284 2176 2322 2240
rect 1702 2160 2322 2176
rect 1702 2096 1740 2160
rect 1804 2096 1820 2160
rect 1884 2096 1900 2160
rect 1964 2096 1980 2160
rect 2044 2096 2060 2160
rect 2124 2096 2140 2160
rect 2204 2096 2220 2160
rect 2284 2096 2322 2160
rect 1702 2080 2322 2096
rect 1702 2016 1740 2080
rect 1804 2016 1820 2080
rect 1884 2016 1900 2080
rect 1964 2016 1980 2080
rect 2044 2016 2060 2080
rect 2124 2016 2140 2080
rect 2204 2016 2220 2080
rect 2284 2016 2322 2080
rect 1702 2000 2322 2016
rect 1702 1936 1740 2000
rect 1804 1936 1820 2000
rect 1884 1936 1900 2000
rect 1964 1936 1980 2000
rect 2044 1936 2060 2000
rect 2124 1936 2140 2000
rect 2204 1936 2220 2000
rect 2284 1936 2322 2000
rect 1702 0 2322 1936
rect 4702 84592 5322 87000
rect 4702 84528 4740 84592
rect 4804 84528 4820 84592
rect 4884 84528 4900 84592
rect 4964 84528 4980 84592
rect 5044 84528 5060 84592
rect 5124 84528 5140 84592
rect 5204 84528 5220 84592
rect 5284 84528 5322 84592
rect 4702 84512 5322 84528
rect 4702 84448 4740 84512
rect 4804 84448 4820 84512
rect 4884 84448 4900 84512
rect 4964 84448 4980 84512
rect 5044 84448 5060 84512
rect 5124 84448 5140 84512
rect 5204 84448 5220 84512
rect 5284 84448 5322 84512
rect 4702 84432 5322 84448
rect 4702 84368 4740 84432
rect 4804 84368 4820 84432
rect 4884 84368 4900 84432
rect 4964 84368 4980 84432
rect 5044 84368 5060 84432
rect 5124 84368 5140 84432
rect 5204 84368 5220 84432
rect 5284 84368 5322 84432
rect 4702 84352 5322 84368
rect 4702 84288 4740 84352
rect 4804 84288 4820 84352
rect 4884 84288 4900 84352
rect 4964 84288 4980 84352
rect 5044 84288 5060 84352
rect 5124 84288 5140 84352
rect 5204 84288 5220 84352
rect 5284 84288 5322 84352
rect 4702 74592 5322 84288
rect 4702 74528 4740 74592
rect 4804 74528 4820 74592
rect 4884 74528 4900 74592
rect 4964 74528 4980 74592
rect 5044 74528 5060 74592
rect 5124 74528 5140 74592
rect 5204 74528 5220 74592
rect 5284 74528 5322 74592
rect 4702 74512 5322 74528
rect 4702 74448 4740 74512
rect 4804 74448 4820 74512
rect 4884 74448 4900 74512
rect 4964 74448 4980 74512
rect 5044 74448 5060 74512
rect 5124 74448 5140 74512
rect 5204 74448 5220 74512
rect 5284 74448 5322 74512
rect 4702 74432 5322 74448
rect 4702 74368 4740 74432
rect 4804 74368 4820 74432
rect 4884 74368 4900 74432
rect 4964 74368 4980 74432
rect 5044 74368 5060 74432
rect 5124 74368 5140 74432
rect 5204 74368 5220 74432
rect 5284 74368 5322 74432
rect 4702 74352 5322 74368
rect 4702 74288 4740 74352
rect 4804 74288 4820 74352
rect 4884 74288 4900 74352
rect 4964 74288 4980 74352
rect 5044 74288 5060 74352
rect 5124 74288 5140 74352
rect 5204 74288 5220 74352
rect 5284 74288 5322 74352
rect 4702 64592 5322 74288
rect 4702 64528 4740 64592
rect 4804 64528 4820 64592
rect 4884 64528 4900 64592
rect 4964 64528 4980 64592
rect 5044 64528 5060 64592
rect 5124 64528 5140 64592
rect 5204 64528 5220 64592
rect 5284 64528 5322 64592
rect 4702 64512 5322 64528
rect 4702 64448 4740 64512
rect 4804 64448 4820 64512
rect 4884 64448 4900 64512
rect 4964 64448 4980 64512
rect 5044 64448 5060 64512
rect 5124 64448 5140 64512
rect 5204 64448 5220 64512
rect 5284 64448 5322 64512
rect 4702 64432 5322 64448
rect 4702 64368 4740 64432
rect 4804 64368 4820 64432
rect 4884 64368 4900 64432
rect 4964 64368 4980 64432
rect 5044 64368 5060 64432
rect 5124 64368 5140 64432
rect 5204 64368 5220 64432
rect 5284 64368 5322 64432
rect 4702 64352 5322 64368
rect 4702 64288 4740 64352
rect 4804 64288 4820 64352
rect 4884 64288 4900 64352
rect 4964 64288 4980 64352
rect 5044 64288 5060 64352
rect 5124 64288 5140 64352
rect 5204 64288 5220 64352
rect 5284 64288 5322 64352
rect 4702 54592 5322 64288
rect 4702 54528 4740 54592
rect 4804 54528 4820 54592
rect 4884 54528 4900 54592
rect 4964 54528 4980 54592
rect 5044 54528 5060 54592
rect 5124 54528 5140 54592
rect 5204 54528 5220 54592
rect 5284 54528 5322 54592
rect 4702 54512 5322 54528
rect 4702 54448 4740 54512
rect 4804 54448 4820 54512
rect 4884 54448 4900 54512
rect 4964 54448 4980 54512
rect 5044 54448 5060 54512
rect 5124 54448 5140 54512
rect 5204 54448 5220 54512
rect 5284 54448 5322 54512
rect 4702 54432 5322 54448
rect 4702 54368 4740 54432
rect 4804 54368 4820 54432
rect 4884 54368 4900 54432
rect 4964 54368 4980 54432
rect 5044 54368 5060 54432
rect 5124 54368 5140 54432
rect 5204 54368 5220 54432
rect 5284 54368 5322 54432
rect 4702 54352 5322 54368
rect 4702 54288 4740 54352
rect 4804 54288 4820 54352
rect 4884 54288 4900 54352
rect 4964 54288 4980 54352
rect 5044 54288 5060 54352
rect 5124 54288 5140 54352
rect 5204 54288 5220 54352
rect 5284 54288 5322 54352
rect 4702 44592 5322 54288
rect 4702 44528 4740 44592
rect 4804 44528 4820 44592
rect 4884 44528 4900 44592
rect 4964 44528 4980 44592
rect 5044 44528 5060 44592
rect 5124 44528 5140 44592
rect 5204 44528 5220 44592
rect 5284 44528 5322 44592
rect 4702 44512 5322 44528
rect 4702 44448 4740 44512
rect 4804 44448 4820 44512
rect 4884 44448 4900 44512
rect 4964 44448 4980 44512
rect 5044 44448 5060 44512
rect 5124 44448 5140 44512
rect 5204 44448 5220 44512
rect 5284 44448 5322 44512
rect 4702 44432 5322 44448
rect 4702 44368 4740 44432
rect 4804 44368 4820 44432
rect 4884 44368 4900 44432
rect 4964 44368 4980 44432
rect 5044 44368 5060 44432
rect 5124 44368 5140 44432
rect 5204 44368 5220 44432
rect 5284 44368 5322 44432
rect 4702 44352 5322 44368
rect 4702 44288 4740 44352
rect 4804 44288 4820 44352
rect 4884 44288 4900 44352
rect 4964 44288 4980 44352
rect 5044 44288 5060 44352
rect 5124 44288 5140 44352
rect 5204 44288 5220 44352
rect 5284 44288 5322 44352
rect 4702 34592 5322 44288
rect 4702 34528 4740 34592
rect 4804 34528 4820 34592
rect 4884 34528 4900 34592
rect 4964 34528 4980 34592
rect 5044 34528 5060 34592
rect 5124 34528 5140 34592
rect 5204 34528 5220 34592
rect 5284 34528 5322 34592
rect 4702 34512 5322 34528
rect 4702 34448 4740 34512
rect 4804 34448 4820 34512
rect 4884 34448 4900 34512
rect 4964 34448 4980 34512
rect 5044 34448 5060 34512
rect 5124 34448 5140 34512
rect 5204 34448 5220 34512
rect 5284 34448 5322 34512
rect 4702 34432 5322 34448
rect 4702 34368 4740 34432
rect 4804 34368 4820 34432
rect 4884 34368 4900 34432
rect 4964 34368 4980 34432
rect 5044 34368 5060 34432
rect 5124 34368 5140 34432
rect 5204 34368 5220 34432
rect 5284 34368 5322 34432
rect 4702 34352 5322 34368
rect 4702 34288 4740 34352
rect 4804 34288 4820 34352
rect 4884 34288 4900 34352
rect 4964 34288 4980 34352
rect 5044 34288 5060 34352
rect 5124 34288 5140 34352
rect 5204 34288 5220 34352
rect 5284 34288 5322 34352
rect 4702 24592 5322 34288
rect 4702 24528 4740 24592
rect 4804 24528 4820 24592
rect 4884 24528 4900 24592
rect 4964 24528 4980 24592
rect 5044 24528 5060 24592
rect 5124 24528 5140 24592
rect 5204 24528 5220 24592
rect 5284 24528 5322 24592
rect 4702 24512 5322 24528
rect 4702 24448 4740 24512
rect 4804 24448 4820 24512
rect 4884 24448 4900 24512
rect 4964 24448 4980 24512
rect 5044 24448 5060 24512
rect 5124 24448 5140 24512
rect 5204 24448 5220 24512
rect 5284 24448 5322 24512
rect 4702 24432 5322 24448
rect 4702 24368 4740 24432
rect 4804 24368 4820 24432
rect 4884 24368 4900 24432
rect 4964 24368 4980 24432
rect 5044 24368 5060 24432
rect 5124 24368 5140 24432
rect 5204 24368 5220 24432
rect 5284 24368 5322 24432
rect 4702 24352 5322 24368
rect 4702 24288 4740 24352
rect 4804 24288 4820 24352
rect 4884 24288 4900 24352
rect 4964 24288 4980 24352
rect 5044 24288 5060 24352
rect 5124 24288 5140 24352
rect 5204 24288 5220 24352
rect 5284 24288 5322 24352
rect 4702 14592 5322 24288
rect 4702 14528 4740 14592
rect 4804 14528 4820 14592
rect 4884 14528 4900 14592
rect 4964 14528 4980 14592
rect 5044 14528 5060 14592
rect 5124 14528 5140 14592
rect 5204 14528 5220 14592
rect 5284 14528 5322 14592
rect 4702 14512 5322 14528
rect 4702 14448 4740 14512
rect 4804 14448 4820 14512
rect 4884 14448 4900 14512
rect 4964 14448 4980 14512
rect 5044 14448 5060 14512
rect 5124 14448 5140 14512
rect 5204 14448 5220 14512
rect 5284 14448 5322 14512
rect 4702 14432 5322 14448
rect 4702 14368 4740 14432
rect 4804 14368 4820 14432
rect 4884 14368 4900 14432
rect 4964 14368 4980 14432
rect 5044 14368 5060 14432
rect 5124 14368 5140 14432
rect 5204 14368 5220 14432
rect 5284 14368 5322 14432
rect 4702 14352 5322 14368
rect 4702 14288 4740 14352
rect 4804 14288 4820 14352
rect 4884 14288 4900 14352
rect 4964 14288 4980 14352
rect 5044 14288 5060 14352
rect 5124 14288 5140 14352
rect 5204 14288 5220 14352
rect 5284 14288 5322 14352
rect 4702 4592 5322 14288
rect 4702 4528 4740 4592
rect 4804 4528 4820 4592
rect 4884 4528 4900 4592
rect 4964 4528 4980 4592
rect 5044 4528 5060 4592
rect 5124 4528 5140 4592
rect 5204 4528 5220 4592
rect 5284 4528 5322 4592
rect 4702 4512 5322 4528
rect 4702 4448 4740 4512
rect 4804 4448 4820 4512
rect 4884 4448 4900 4512
rect 4964 4448 4980 4512
rect 5044 4448 5060 4512
rect 5124 4448 5140 4512
rect 5204 4448 5220 4512
rect 5284 4448 5322 4512
rect 4702 4432 5322 4448
rect 4702 4368 4740 4432
rect 4804 4368 4820 4432
rect 4884 4368 4900 4432
rect 4964 4368 4980 4432
rect 5044 4368 5060 4432
rect 5124 4368 5140 4432
rect 5204 4368 5220 4432
rect 5284 4368 5322 4432
rect 4702 4352 5322 4368
rect 4702 4288 4740 4352
rect 4804 4288 4820 4352
rect 4884 4288 4900 4352
rect 4964 4288 4980 4352
rect 5044 4288 5060 4352
rect 5124 4288 5140 4352
rect 5204 4288 5220 4352
rect 5284 4288 5322 4352
rect 4702 0 5322 4288
rect 7702 82240 8322 87000
rect 7702 82176 7740 82240
rect 7804 82176 7820 82240
rect 7884 82176 7900 82240
rect 7964 82176 7980 82240
rect 8044 82176 8060 82240
rect 8124 82176 8140 82240
rect 8204 82176 8220 82240
rect 8284 82176 8322 82240
rect 7702 82160 8322 82176
rect 7702 82096 7740 82160
rect 7804 82096 7820 82160
rect 7884 82096 7900 82160
rect 7964 82096 7980 82160
rect 8044 82096 8060 82160
rect 8124 82096 8140 82160
rect 8204 82096 8220 82160
rect 8284 82096 8322 82160
rect 7702 82080 8322 82096
rect 7702 82016 7740 82080
rect 7804 82016 7820 82080
rect 7884 82016 7900 82080
rect 7964 82016 7980 82080
rect 8044 82016 8060 82080
rect 8124 82016 8140 82080
rect 8204 82016 8220 82080
rect 8284 82016 8322 82080
rect 7702 82000 8322 82016
rect 7702 81936 7740 82000
rect 7804 81936 7820 82000
rect 7884 81936 7900 82000
rect 7964 81936 7980 82000
rect 8044 81936 8060 82000
rect 8124 81936 8140 82000
rect 8204 81936 8220 82000
rect 8284 81936 8322 82000
rect 7702 72240 8322 81936
rect 7702 72176 7740 72240
rect 7804 72176 7820 72240
rect 7884 72176 7900 72240
rect 7964 72176 7980 72240
rect 8044 72176 8060 72240
rect 8124 72176 8140 72240
rect 8204 72176 8220 72240
rect 8284 72176 8322 72240
rect 7702 72160 8322 72176
rect 7702 72096 7740 72160
rect 7804 72096 7820 72160
rect 7884 72096 7900 72160
rect 7964 72096 7980 72160
rect 8044 72096 8060 72160
rect 8124 72096 8140 72160
rect 8204 72096 8220 72160
rect 8284 72096 8322 72160
rect 7702 72080 8322 72096
rect 7702 72016 7740 72080
rect 7804 72016 7820 72080
rect 7884 72016 7900 72080
rect 7964 72016 7980 72080
rect 8044 72016 8060 72080
rect 8124 72016 8140 72080
rect 8204 72016 8220 72080
rect 8284 72016 8322 72080
rect 7702 72000 8322 72016
rect 7702 71936 7740 72000
rect 7804 71936 7820 72000
rect 7884 71936 7900 72000
rect 7964 71936 7980 72000
rect 8044 71936 8060 72000
rect 8124 71936 8140 72000
rect 8204 71936 8220 72000
rect 8284 71936 8322 72000
rect 7702 62240 8322 71936
rect 7702 62176 7740 62240
rect 7804 62176 7820 62240
rect 7884 62176 7900 62240
rect 7964 62176 7980 62240
rect 8044 62176 8060 62240
rect 8124 62176 8140 62240
rect 8204 62176 8220 62240
rect 8284 62176 8322 62240
rect 7702 62160 8322 62176
rect 7702 62096 7740 62160
rect 7804 62096 7820 62160
rect 7884 62096 7900 62160
rect 7964 62096 7980 62160
rect 8044 62096 8060 62160
rect 8124 62096 8140 62160
rect 8204 62096 8220 62160
rect 8284 62096 8322 62160
rect 7702 62080 8322 62096
rect 7702 62016 7740 62080
rect 7804 62016 7820 62080
rect 7884 62016 7900 62080
rect 7964 62016 7980 62080
rect 8044 62016 8060 62080
rect 8124 62016 8140 62080
rect 8204 62016 8220 62080
rect 8284 62016 8322 62080
rect 7702 62000 8322 62016
rect 7702 61936 7740 62000
rect 7804 61936 7820 62000
rect 7884 61936 7900 62000
rect 7964 61936 7980 62000
rect 8044 61936 8060 62000
rect 8124 61936 8140 62000
rect 8204 61936 8220 62000
rect 8284 61936 8322 62000
rect 7702 52240 8322 61936
rect 7702 52176 7740 52240
rect 7804 52176 7820 52240
rect 7884 52176 7900 52240
rect 7964 52176 7980 52240
rect 8044 52176 8060 52240
rect 8124 52176 8140 52240
rect 8204 52176 8220 52240
rect 8284 52176 8322 52240
rect 7702 52160 8322 52176
rect 7702 52096 7740 52160
rect 7804 52096 7820 52160
rect 7884 52096 7900 52160
rect 7964 52096 7980 52160
rect 8044 52096 8060 52160
rect 8124 52096 8140 52160
rect 8204 52096 8220 52160
rect 8284 52096 8322 52160
rect 7702 52080 8322 52096
rect 7702 52016 7740 52080
rect 7804 52016 7820 52080
rect 7884 52016 7900 52080
rect 7964 52016 7980 52080
rect 8044 52016 8060 52080
rect 8124 52016 8140 52080
rect 8204 52016 8220 52080
rect 8284 52016 8322 52080
rect 7702 52000 8322 52016
rect 7702 51936 7740 52000
rect 7804 51936 7820 52000
rect 7884 51936 7900 52000
rect 7964 51936 7980 52000
rect 8044 51936 8060 52000
rect 8124 51936 8140 52000
rect 8204 51936 8220 52000
rect 8284 51936 8322 52000
rect 7702 42240 8322 51936
rect 7702 42176 7740 42240
rect 7804 42176 7820 42240
rect 7884 42176 7900 42240
rect 7964 42176 7980 42240
rect 8044 42176 8060 42240
rect 8124 42176 8140 42240
rect 8204 42176 8220 42240
rect 8284 42176 8322 42240
rect 7702 42160 8322 42176
rect 7702 42096 7740 42160
rect 7804 42096 7820 42160
rect 7884 42096 7900 42160
rect 7964 42096 7980 42160
rect 8044 42096 8060 42160
rect 8124 42096 8140 42160
rect 8204 42096 8220 42160
rect 8284 42096 8322 42160
rect 7702 42080 8322 42096
rect 7702 42016 7740 42080
rect 7804 42016 7820 42080
rect 7884 42016 7900 42080
rect 7964 42016 7980 42080
rect 8044 42016 8060 42080
rect 8124 42016 8140 42080
rect 8204 42016 8220 42080
rect 8284 42016 8322 42080
rect 7702 42000 8322 42016
rect 7702 41936 7740 42000
rect 7804 41936 7820 42000
rect 7884 41936 7900 42000
rect 7964 41936 7980 42000
rect 8044 41936 8060 42000
rect 8124 41936 8140 42000
rect 8204 41936 8220 42000
rect 8284 41936 8322 42000
rect 7702 32240 8322 41936
rect 7702 32176 7740 32240
rect 7804 32176 7820 32240
rect 7884 32176 7900 32240
rect 7964 32176 7980 32240
rect 8044 32176 8060 32240
rect 8124 32176 8140 32240
rect 8204 32176 8220 32240
rect 8284 32176 8322 32240
rect 7702 32160 8322 32176
rect 7702 32096 7740 32160
rect 7804 32096 7820 32160
rect 7884 32096 7900 32160
rect 7964 32096 7980 32160
rect 8044 32096 8060 32160
rect 8124 32096 8140 32160
rect 8204 32096 8220 32160
rect 8284 32096 8322 32160
rect 7702 32080 8322 32096
rect 7702 32016 7740 32080
rect 7804 32016 7820 32080
rect 7884 32016 7900 32080
rect 7964 32016 7980 32080
rect 8044 32016 8060 32080
rect 8124 32016 8140 32080
rect 8204 32016 8220 32080
rect 8284 32016 8322 32080
rect 7702 32000 8322 32016
rect 7702 31936 7740 32000
rect 7804 31936 7820 32000
rect 7884 31936 7900 32000
rect 7964 31936 7980 32000
rect 8044 31936 8060 32000
rect 8124 31936 8140 32000
rect 8204 31936 8220 32000
rect 8284 31936 8322 32000
rect 7702 22240 8322 31936
rect 7702 22176 7740 22240
rect 7804 22176 7820 22240
rect 7884 22176 7900 22240
rect 7964 22176 7980 22240
rect 8044 22176 8060 22240
rect 8124 22176 8140 22240
rect 8204 22176 8220 22240
rect 8284 22176 8322 22240
rect 7702 22160 8322 22176
rect 7702 22096 7740 22160
rect 7804 22096 7820 22160
rect 7884 22096 7900 22160
rect 7964 22096 7980 22160
rect 8044 22096 8060 22160
rect 8124 22096 8140 22160
rect 8204 22096 8220 22160
rect 8284 22096 8322 22160
rect 7702 22080 8322 22096
rect 7702 22016 7740 22080
rect 7804 22016 7820 22080
rect 7884 22016 7900 22080
rect 7964 22016 7980 22080
rect 8044 22016 8060 22080
rect 8124 22016 8140 22080
rect 8204 22016 8220 22080
rect 8284 22016 8322 22080
rect 7702 22000 8322 22016
rect 7702 21936 7740 22000
rect 7804 21936 7820 22000
rect 7884 21936 7900 22000
rect 7964 21936 7980 22000
rect 8044 21936 8060 22000
rect 8124 21936 8140 22000
rect 8204 21936 8220 22000
rect 8284 21936 8322 22000
rect 7702 12240 8322 21936
rect 7702 12176 7740 12240
rect 7804 12176 7820 12240
rect 7884 12176 7900 12240
rect 7964 12176 7980 12240
rect 8044 12176 8060 12240
rect 8124 12176 8140 12240
rect 8204 12176 8220 12240
rect 8284 12176 8322 12240
rect 7702 12160 8322 12176
rect 7702 12096 7740 12160
rect 7804 12096 7820 12160
rect 7884 12096 7900 12160
rect 7964 12096 7980 12160
rect 8044 12096 8060 12160
rect 8124 12096 8140 12160
rect 8204 12096 8220 12160
rect 8284 12096 8322 12160
rect 7702 12080 8322 12096
rect 7702 12016 7740 12080
rect 7804 12016 7820 12080
rect 7884 12016 7900 12080
rect 7964 12016 7980 12080
rect 8044 12016 8060 12080
rect 8124 12016 8140 12080
rect 8204 12016 8220 12080
rect 8284 12016 8322 12080
rect 7702 12000 8322 12016
rect 7702 11936 7740 12000
rect 7804 11936 7820 12000
rect 7884 11936 7900 12000
rect 7964 11936 7980 12000
rect 8044 11936 8060 12000
rect 8124 11936 8140 12000
rect 8204 11936 8220 12000
rect 8284 11936 8322 12000
rect 7702 2240 8322 11936
rect 7702 2176 7740 2240
rect 7804 2176 7820 2240
rect 7884 2176 7900 2240
rect 7964 2176 7980 2240
rect 8044 2176 8060 2240
rect 8124 2176 8140 2240
rect 8204 2176 8220 2240
rect 8284 2176 8322 2240
rect 7702 2160 8322 2176
rect 7702 2096 7740 2160
rect 7804 2096 7820 2160
rect 7884 2096 7900 2160
rect 7964 2096 7980 2160
rect 8044 2096 8060 2160
rect 8124 2096 8140 2160
rect 8204 2096 8220 2160
rect 8284 2096 8322 2160
rect 7702 2080 8322 2096
rect 7702 2016 7740 2080
rect 7804 2016 7820 2080
rect 7884 2016 7900 2080
rect 7964 2016 7980 2080
rect 8044 2016 8060 2080
rect 8124 2016 8140 2080
rect 8204 2016 8220 2080
rect 8284 2016 8322 2080
rect 7702 2000 8322 2016
rect 7702 1936 7740 2000
rect 7804 1936 7820 2000
rect 7884 1936 7900 2000
rect 7964 1936 7980 2000
rect 8044 1936 8060 2000
rect 8124 1936 8140 2000
rect 8204 1936 8220 2000
rect 8284 1936 8322 2000
rect 7702 0 8322 1936
rect 10702 84592 11322 87000
rect 10702 84528 10740 84592
rect 10804 84528 10820 84592
rect 10884 84528 10900 84592
rect 10964 84528 10980 84592
rect 11044 84528 11060 84592
rect 11124 84528 11140 84592
rect 11204 84528 11220 84592
rect 11284 84528 11322 84592
rect 10702 84512 11322 84528
rect 10702 84448 10740 84512
rect 10804 84448 10820 84512
rect 10884 84448 10900 84512
rect 10964 84448 10980 84512
rect 11044 84448 11060 84512
rect 11124 84448 11140 84512
rect 11204 84448 11220 84512
rect 11284 84448 11322 84512
rect 10702 84432 11322 84448
rect 10702 84368 10740 84432
rect 10804 84368 10820 84432
rect 10884 84368 10900 84432
rect 10964 84368 10980 84432
rect 11044 84368 11060 84432
rect 11124 84368 11140 84432
rect 11204 84368 11220 84432
rect 11284 84368 11322 84432
rect 10702 84352 11322 84368
rect 10702 84288 10740 84352
rect 10804 84288 10820 84352
rect 10884 84288 10900 84352
rect 10964 84288 10980 84352
rect 11044 84288 11060 84352
rect 11124 84288 11140 84352
rect 11204 84288 11220 84352
rect 11284 84288 11322 84352
rect 10702 74592 11322 84288
rect 10702 74528 10740 74592
rect 10804 74528 10820 74592
rect 10884 74528 10900 74592
rect 10964 74528 10980 74592
rect 11044 74528 11060 74592
rect 11124 74528 11140 74592
rect 11204 74528 11220 74592
rect 11284 74528 11322 74592
rect 10702 74512 11322 74528
rect 10702 74448 10740 74512
rect 10804 74448 10820 74512
rect 10884 74448 10900 74512
rect 10964 74448 10980 74512
rect 11044 74448 11060 74512
rect 11124 74448 11140 74512
rect 11204 74448 11220 74512
rect 11284 74448 11322 74512
rect 10702 74432 11322 74448
rect 10702 74368 10740 74432
rect 10804 74368 10820 74432
rect 10884 74368 10900 74432
rect 10964 74368 10980 74432
rect 11044 74368 11060 74432
rect 11124 74368 11140 74432
rect 11204 74368 11220 74432
rect 11284 74368 11322 74432
rect 10702 74352 11322 74368
rect 10702 74288 10740 74352
rect 10804 74288 10820 74352
rect 10884 74288 10900 74352
rect 10964 74288 10980 74352
rect 11044 74288 11060 74352
rect 11124 74288 11140 74352
rect 11204 74288 11220 74352
rect 11284 74288 11322 74352
rect 10702 64592 11322 74288
rect 10702 64528 10740 64592
rect 10804 64528 10820 64592
rect 10884 64528 10900 64592
rect 10964 64528 10980 64592
rect 11044 64528 11060 64592
rect 11124 64528 11140 64592
rect 11204 64528 11220 64592
rect 11284 64528 11322 64592
rect 10702 64512 11322 64528
rect 10702 64448 10740 64512
rect 10804 64448 10820 64512
rect 10884 64448 10900 64512
rect 10964 64448 10980 64512
rect 11044 64448 11060 64512
rect 11124 64448 11140 64512
rect 11204 64448 11220 64512
rect 11284 64448 11322 64512
rect 10702 64432 11322 64448
rect 10702 64368 10740 64432
rect 10804 64368 10820 64432
rect 10884 64368 10900 64432
rect 10964 64368 10980 64432
rect 11044 64368 11060 64432
rect 11124 64368 11140 64432
rect 11204 64368 11220 64432
rect 11284 64368 11322 64432
rect 10702 64352 11322 64368
rect 10702 64288 10740 64352
rect 10804 64288 10820 64352
rect 10884 64288 10900 64352
rect 10964 64288 10980 64352
rect 11044 64288 11060 64352
rect 11124 64288 11140 64352
rect 11204 64288 11220 64352
rect 11284 64288 11322 64352
rect 10702 54592 11322 64288
rect 10702 54528 10740 54592
rect 10804 54528 10820 54592
rect 10884 54528 10900 54592
rect 10964 54528 10980 54592
rect 11044 54528 11060 54592
rect 11124 54528 11140 54592
rect 11204 54528 11220 54592
rect 11284 54528 11322 54592
rect 10702 54512 11322 54528
rect 10702 54448 10740 54512
rect 10804 54448 10820 54512
rect 10884 54448 10900 54512
rect 10964 54448 10980 54512
rect 11044 54448 11060 54512
rect 11124 54448 11140 54512
rect 11204 54448 11220 54512
rect 11284 54448 11322 54512
rect 10702 54432 11322 54448
rect 10702 54368 10740 54432
rect 10804 54368 10820 54432
rect 10884 54368 10900 54432
rect 10964 54368 10980 54432
rect 11044 54368 11060 54432
rect 11124 54368 11140 54432
rect 11204 54368 11220 54432
rect 11284 54368 11322 54432
rect 10702 54352 11322 54368
rect 10702 54288 10740 54352
rect 10804 54288 10820 54352
rect 10884 54288 10900 54352
rect 10964 54288 10980 54352
rect 11044 54288 11060 54352
rect 11124 54288 11140 54352
rect 11204 54288 11220 54352
rect 11284 54288 11322 54352
rect 10702 44592 11322 54288
rect 10702 44528 10740 44592
rect 10804 44528 10820 44592
rect 10884 44528 10900 44592
rect 10964 44528 10980 44592
rect 11044 44528 11060 44592
rect 11124 44528 11140 44592
rect 11204 44528 11220 44592
rect 11284 44528 11322 44592
rect 10702 44512 11322 44528
rect 10702 44448 10740 44512
rect 10804 44448 10820 44512
rect 10884 44448 10900 44512
rect 10964 44448 10980 44512
rect 11044 44448 11060 44512
rect 11124 44448 11140 44512
rect 11204 44448 11220 44512
rect 11284 44448 11322 44512
rect 10702 44432 11322 44448
rect 10702 44368 10740 44432
rect 10804 44368 10820 44432
rect 10884 44368 10900 44432
rect 10964 44368 10980 44432
rect 11044 44368 11060 44432
rect 11124 44368 11140 44432
rect 11204 44368 11220 44432
rect 11284 44368 11322 44432
rect 10702 44352 11322 44368
rect 10702 44288 10740 44352
rect 10804 44288 10820 44352
rect 10884 44288 10900 44352
rect 10964 44288 10980 44352
rect 11044 44288 11060 44352
rect 11124 44288 11140 44352
rect 11204 44288 11220 44352
rect 11284 44288 11322 44352
rect 10702 34592 11322 44288
rect 10702 34528 10740 34592
rect 10804 34528 10820 34592
rect 10884 34528 10900 34592
rect 10964 34528 10980 34592
rect 11044 34528 11060 34592
rect 11124 34528 11140 34592
rect 11204 34528 11220 34592
rect 11284 34528 11322 34592
rect 10702 34512 11322 34528
rect 10702 34448 10740 34512
rect 10804 34448 10820 34512
rect 10884 34448 10900 34512
rect 10964 34448 10980 34512
rect 11044 34448 11060 34512
rect 11124 34448 11140 34512
rect 11204 34448 11220 34512
rect 11284 34448 11322 34512
rect 10702 34432 11322 34448
rect 10702 34368 10740 34432
rect 10804 34368 10820 34432
rect 10884 34368 10900 34432
rect 10964 34368 10980 34432
rect 11044 34368 11060 34432
rect 11124 34368 11140 34432
rect 11204 34368 11220 34432
rect 11284 34368 11322 34432
rect 10702 34352 11322 34368
rect 10702 34288 10740 34352
rect 10804 34288 10820 34352
rect 10884 34288 10900 34352
rect 10964 34288 10980 34352
rect 11044 34288 11060 34352
rect 11124 34288 11140 34352
rect 11204 34288 11220 34352
rect 11284 34288 11322 34352
rect 10702 24592 11322 34288
rect 10702 24528 10740 24592
rect 10804 24528 10820 24592
rect 10884 24528 10900 24592
rect 10964 24528 10980 24592
rect 11044 24528 11060 24592
rect 11124 24528 11140 24592
rect 11204 24528 11220 24592
rect 11284 24528 11322 24592
rect 10702 24512 11322 24528
rect 10702 24448 10740 24512
rect 10804 24448 10820 24512
rect 10884 24448 10900 24512
rect 10964 24448 10980 24512
rect 11044 24448 11060 24512
rect 11124 24448 11140 24512
rect 11204 24448 11220 24512
rect 11284 24448 11322 24512
rect 10702 24432 11322 24448
rect 10702 24368 10740 24432
rect 10804 24368 10820 24432
rect 10884 24368 10900 24432
rect 10964 24368 10980 24432
rect 11044 24368 11060 24432
rect 11124 24368 11140 24432
rect 11204 24368 11220 24432
rect 11284 24368 11322 24432
rect 10702 24352 11322 24368
rect 10702 24288 10740 24352
rect 10804 24288 10820 24352
rect 10884 24288 10900 24352
rect 10964 24288 10980 24352
rect 11044 24288 11060 24352
rect 11124 24288 11140 24352
rect 11204 24288 11220 24352
rect 11284 24288 11322 24352
rect 10702 14592 11322 24288
rect 10702 14528 10740 14592
rect 10804 14528 10820 14592
rect 10884 14528 10900 14592
rect 10964 14528 10980 14592
rect 11044 14528 11060 14592
rect 11124 14528 11140 14592
rect 11204 14528 11220 14592
rect 11284 14528 11322 14592
rect 10702 14512 11322 14528
rect 10702 14448 10740 14512
rect 10804 14448 10820 14512
rect 10884 14448 10900 14512
rect 10964 14448 10980 14512
rect 11044 14448 11060 14512
rect 11124 14448 11140 14512
rect 11204 14448 11220 14512
rect 11284 14448 11322 14512
rect 10702 14432 11322 14448
rect 10702 14368 10740 14432
rect 10804 14368 10820 14432
rect 10884 14368 10900 14432
rect 10964 14368 10980 14432
rect 11044 14368 11060 14432
rect 11124 14368 11140 14432
rect 11204 14368 11220 14432
rect 11284 14368 11322 14432
rect 10702 14352 11322 14368
rect 10702 14288 10740 14352
rect 10804 14288 10820 14352
rect 10884 14288 10900 14352
rect 10964 14288 10980 14352
rect 11044 14288 11060 14352
rect 11124 14288 11140 14352
rect 11204 14288 11220 14352
rect 11284 14288 11322 14352
rect 10702 4592 11322 14288
rect 10702 4528 10740 4592
rect 10804 4528 10820 4592
rect 10884 4528 10900 4592
rect 10964 4528 10980 4592
rect 11044 4528 11060 4592
rect 11124 4528 11140 4592
rect 11204 4528 11220 4592
rect 11284 4528 11322 4592
rect 10702 4512 11322 4528
rect 10702 4448 10740 4512
rect 10804 4448 10820 4512
rect 10884 4448 10900 4512
rect 10964 4448 10980 4512
rect 11044 4448 11060 4512
rect 11124 4448 11140 4512
rect 11204 4448 11220 4512
rect 11284 4448 11322 4512
rect 10702 4432 11322 4448
rect 10702 4368 10740 4432
rect 10804 4368 10820 4432
rect 10884 4368 10900 4432
rect 10964 4368 10980 4432
rect 11044 4368 11060 4432
rect 11124 4368 11140 4432
rect 11204 4368 11220 4432
rect 11284 4368 11322 4432
rect 10702 4352 11322 4368
rect 10702 4288 10740 4352
rect 10804 4288 10820 4352
rect 10884 4288 10900 4352
rect 10964 4288 10980 4352
rect 11044 4288 11060 4352
rect 11124 4288 11140 4352
rect 11204 4288 11220 4352
rect 11284 4288 11322 4352
rect 10702 0 11322 4288
rect 13702 82240 14322 87000
rect 13702 82176 13740 82240
rect 13804 82176 13820 82240
rect 13884 82176 13900 82240
rect 13964 82176 13980 82240
rect 14044 82176 14060 82240
rect 14124 82176 14140 82240
rect 14204 82176 14220 82240
rect 14284 82176 14322 82240
rect 13702 82160 14322 82176
rect 13702 82096 13740 82160
rect 13804 82096 13820 82160
rect 13884 82096 13900 82160
rect 13964 82096 13980 82160
rect 14044 82096 14060 82160
rect 14124 82096 14140 82160
rect 14204 82096 14220 82160
rect 14284 82096 14322 82160
rect 13702 82080 14322 82096
rect 13702 82016 13740 82080
rect 13804 82016 13820 82080
rect 13884 82016 13900 82080
rect 13964 82016 13980 82080
rect 14044 82016 14060 82080
rect 14124 82016 14140 82080
rect 14204 82016 14220 82080
rect 14284 82016 14322 82080
rect 13702 82000 14322 82016
rect 13702 81936 13740 82000
rect 13804 81936 13820 82000
rect 13884 81936 13900 82000
rect 13964 81936 13980 82000
rect 14044 81936 14060 82000
rect 14124 81936 14140 82000
rect 14204 81936 14220 82000
rect 14284 81936 14322 82000
rect 13702 72240 14322 81936
rect 13702 72176 13740 72240
rect 13804 72176 13820 72240
rect 13884 72176 13900 72240
rect 13964 72176 13980 72240
rect 14044 72176 14060 72240
rect 14124 72176 14140 72240
rect 14204 72176 14220 72240
rect 14284 72176 14322 72240
rect 13702 72160 14322 72176
rect 13702 72096 13740 72160
rect 13804 72096 13820 72160
rect 13884 72096 13900 72160
rect 13964 72096 13980 72160
rect 14044 72096 14060 72160
rect 14124 72096 14140 72160
rect 14204 72096 14220 72160
rect 14284 72096 14322 72160
rect 13702 72080 14322 72096
rect 13702 72016 13740 72080
rect 13804 72016 13820 72080
rect 13884 72016 13900 72080
rect 13964 72016 13980 72080
rect 14044 72016 14060 72080
rect 14124 72016 14140 72080
rect 14204 72016 14220 72080
rect 14284 72016 14322 72080
rect 13702 72000 14322 72016
rect 13702 71936 13740 72000
rect 13804 71936 13820 72000
rect 13884 71936 13900 72000
rect 13964 71936 13980 72000
rect 14044 71936 14060 72000
rect 14124 71936 14140 72000
rect 14204 71936 14220 72000
rect 14284 71936 14322 72000
rect 13702 62240 14322 71936
rect 13702 62176 13740 62240
rect 13804 62176 13820 62240
rect 13884 62176 13900 62240
rect 13964 62176 13980 62240
rect 14044 62176 14060 62240
rect 14124 62176 14140 62240
rect 14204 62176 14220 62240
rect 14284 62176 14322 62240
rect 13702 62160 14322 62176
rect 13702 62096 13740 62160
rect 13804 62096 13820 62160
rect 13884 62096 13900 62160
rect 13964 62096 13980 62160
rect 14044 62096 14060 62160
rect 14124 62096 14140 62160
rect 14204 62096 14220 62160
rect 14284 62096 14322 62160
rect 13702 62080 14322 62096
rect 13702 62016 13740 62080
rect 13804 62016 13820 62080
rect 13884 62016 13900 62080
rect 13964 62016 13980 62080
rect 14044 62016 14060 62080
rect 14124 62016 14140 62080
rect 14204 62016 14220 62080
rect 14284 62016 14322 62080
rect 13702 62000 14322 62016
rect 13702 61936 13740 62000
rect 13804 61936 13820 62000
rect 13884 61936 13900 62000
rect 13964 61936 13980 62000
rect 14044 61936 14060 62000
rect 14124 61936 14140 62000
rect 14204 61936 14220 62000
rect 14284 61936 14322 62000
rect 13702 52240 14322 61936
rect 13702 52176 13740 52240
rect 13804 52176 13820 52240
rect 13884 52176 13900 52240
rect 13964 52176 13980 52240
rect 14044 52176 14060 52240
rect 14124 52176 14140 52240
rect 14204 52176 14220 52240
rect 14284 52176 14322 52240
rect 13702 52160 14322 52176
rect 13702 52096 13740 52160
rect 13804 52096 13820 52160
rect 13884 52096 13900 52160
rect 13964 52096 13980 52160
rect 14044 52096 14060 52160
rect 14124 52096 14140 52160
rect 14204 52096 14220 52160
rect 14284 52096 14322 52160
rect 13702 52080 14322 52096
rect 13702 52016 13740 52080
rect 13804 52016 13820 52080
rect 13884 52016 13900 52080
rect 13964 52016 13980 52080
rect 14044 52016 14060 52080
rect 14124 52016 14140 52080
rect 14204 52016 14220 52080
rect 14284 52016 14322 52080
rect 13702 52000 14322 52016
rect 13702 51936 13740 52000
rect 13804 51936 13820 52000
rect 13884 51936 13900 52000
rect 13964 51936 13980 52000
rect 14044 51936 14060 52000
rect 14124 51936 14140 52000
rect 14204 51936 14220 52000
rect 14284 51936 14322 52000
rect 13702 42240 14322 51936
rect 13702 42176 13740 42240
rect 13804 42176 13820 42240
rect 13884 42176 13900 42240
rect 13964 42176 13980 42240
rect 14044 42176 14060 42240
rect 14124 42176 14140 42240
rect 14204 42176 14220 42240
rect 14284 42176 14322 42240
rect 13702 42160 14322 42176
rect 13702 42096 13740 42160
rect 13804 42096 13820 42160
rect 13884 42096 13900 42160
rect 13964 42096 13980 42160
rect 14044 42096 14060 42160
rect 14124 42096 14140 42160
rect 14204 42096 14220 42160
rect 14284 42096 14322 42160
rect 13702 42080 14322 42096
rect 13702 42016 13740 42080
rect 13804 42016 13820 42080
rect 13884 42016 13900 42080
rect 13964 42016 13980 42080
rect 14044 42016 14060 42080
rect 14124 42016 14140 42080
rect 14204 42016 14220 42080
rect 14284 42016 14322 42080
rect 13702 42000 14322 42016
rect 13702 41936 13740 42000
rect 13804 41936 13820 42000
rect 13884 41936 13900 42000
rect 13964 41936 13980 42000
rect 14044 41936 14060 42000
rect 14124 41936 14140 42000
rect 14204 41936 14220 42000
rect 14284 41936 14322 42000
rect 13702 32240 14322 41936
rect 13702 32176 13740 32240
rect 13804 32176 13820 32240
rect 13884 32176 13900 32240
rect 13964 32176 13980 32240
rect 14044 32176 14060 32240
rect 14124 32176 14140 32240
rect 14204 32176 14220 32240
rect 14284 32176 14322 32240
rect 13702 32160 14322 32176
rect 13702 32096 13740 32160
rect 13804 32096 13820 32160
rect 13884 32096 13900 32160
rect 13964 32096 13980 32160
rect 14044 32096 14060 32160
rect 14124 32096 14140 32160
rect 14204 32096 14220 32160
rect 14284 32096 14322 32160
rect 13702 32080 14322 32096
rect 13702 32016 13740 32080
rect 13804 32016 13820 32080
rect 13884 32016 13900 32080
rect 13964 32016 13980 32080
rect 14044 32016 14060 32080
rect 14124 32016 14140 32080
rect 14204 32016 14220 32080
rect 14284 32016 14322 32080
rect 13702 32000 14322 32016
rect 13702 31936 13740 32000
rect 13804 31936 13820 32000
rect 13884 31936 13900 32000
rect 13964 31936 13980 32000
rect 14044 31936 14060 32000
rect 14124 31936 14140 32000
rect 14204 31936 14220 32000
rect 14284 31936 14322 32000
rect 13702 22240 14322 31936
rect 13702 22176 13740 22240
rect 13804 22176 13820 22240
rect 13884 22176 13900 22240
rect 13964 22176 13980 22240
rect 14044 22176 14060 22240
rect 14124 22176 14140 22240
rect 14204 22176 14220 22240
rect 14284 22176 14322 22240
rect 13702 22160 14322 22176
rect 13702 22096 13740 22160
rect 13804 22096 13820 22160
rect 13884 22096 13900 22160
rect 13964 22096 13980 22160
rect 14044 22096 14060 22160
rect 14124 22096 14140 22160
rect 14204 22096 14220 22160
rect 14284 22096 14322 22160
rect 13702 22080 14322 22096
rect 13702 22016 13740 22080
rect 13804 22016 13820 22080
rect 13884 22016 13900 22080
rect 13964 22016 13980 22080
rect 14044 22016 14060 22080
rect 14124 22016 14140 22080
rect 14204 22016 14220 22080
rect 14284 22016 14322 22080
rect 13702 22000 14322 22016
rect 13702 21936 13740 22000
rect 13804 21936 13820 22000
rect 13884 21936 13900 22000
rect 13964 21936 13980 22000
rect 14044 21936 14060 22000
rect 14124 21936 14140 22000
rect 14204 21936 14220 22000
rect 14284 21936 14322 22000
rect 13702 12240 14322 21936
rect 13702 12176 13740 12240
rect 13804 12176 13820 12240
rect 13884 12176 13900 12240
rect 13964 12176 13980 12240
rect 14044 12176 14060 12240
rect 14124 12176 14140 12240
rect 14204 12176 14220 12240
rect 14284 12176 14322 12240
rect 13702 12160 14322 12176
rect 13702 12096 13740 12160
rect 13804 12096 13820 12160
rect 13884 12096 13900 12160
rect 13964 12096 13980 12160
rect 14044 12096 14060 12160
rect 14124 12096 14140 12160
rect 14204 12096 14220 12160
rect 14284 12096 14322 12160
rect 13702 12080 14322 12096
rect 13702 12016 13740 12080
rect 13804 12016 13820 12080
rect 13884 12016 13900 12080
rect 13964 12016 13980 12080
rect 14044 12016 14060 12080
rect 14124 12016 14140 12080
rect 14204 12016 14220 12080
rect 14284 12016 14322 12080
rect 13702 12000 14322 12016
rect 13702 11936 13740 12000
rect 13804 11936 13820 12000
rect 13884 11936 13900 12000
rect 13964 11936 13980 12000
rect 14044 11936 14060 12000
rect 14124 11936 14140 12000
rect 14204 11936 14220 12000
rect 14284 11936 14322 12000
rect 13702 2240 14322 11936
rect 13702 2176 13740 2240
rect 13804 2176 13820 2240
rect 13884 2176 13900 2240
rect 13964 2176 13980 2240
rect 14044 2176 14060 2240
rect 14124 2176 14140 2240
rect 14204 2176 14220 2240
rect 14284 2176 14322 2240
rect 13702 2160 14322 2176
rect 13702 2096 13740 2160
rect 13804 2096 13820 2160
rect 13884 2096 13900 2160
rect 13964 2096 13980 2160
rect 14044 2096 14060 2160
rect 14124 2096 14140 2160
rect 14204 2096 14220 2160
rect 14284 2096 14322 2160
rect 13702 2080 14322 2096
rect 13702 2016 13740 2080
rect 13804 2016 13820 2080
rect 13884 2016 13900 2080
rect 13964 2016 13980 2080
rect 14044 2016 14060 2080
rect 14124 2016 14140 2080
rect 14204 2016 14220 2080
rect 14284 2016 14322 2080
rect 13702 2000 14322 2016
rect 13702 1936 13740 2000
rect 13804 1936 13820 2000
rect 13884 1936 13900 2000
rect 13964 1936 13980 2000
rect 14044 1936 14060 2000
rect 14124 1936 14140 2000
rect 14204 1936 14220 2000
rect 14284 1936 14322 2000
rect 13702 0 14322 1936
rect 16702 84592 17322 87000
rect 16702 84528 16740 84592
rect 16804 84528 16820 84592
rect 16884 84528 16900 84592
rect 16964 84528 16980 84592
rect 17044 84528 17060 84592
rect 17124 84528 17140 84592
rect 17204 84528 17220 84592
rect 17284 84528 17322 84592
rect 16702 84512 17322 84528
rect 16702 84448 16740 84512
rect 16804 84448 16820 84512
rect 16884 84448 16900 84512
rect 16964 84448 16980 84512
rect 17044 84448 17060 84512
rect 17124 84448 17140 84512
rect 17204 84448 17220 84512
rect 17284 84448 17322 84512
rect 16702 84432 17322 84448
rect 16702 84368 16740 84432
rect 16804 84368 16820 84432
rect 16884 84368 16900 84432
rect 16964 84368 16980 84432
rect 17044 84368 17060 84432
rect 17124 84368 17140 84432
rect 17204 84368 17220 84432
rect 17284 84368 17322 84432
rect 16702 84352 17322 84368
rect 16702 84288 16740 84352
rect 16804 84288 16820 84352
rect 16884 84288 16900 84352
rect 16964 84288 16980 84352
rect 17044 84288 17060 84352
rect 17124 84288 17140 84352
rect 17204 84288 17220 84352
rect 17284 84288 17322 84352
rect 16702 74592 17322 84288
rect 16702 74528 16740 74592
rect 16804 74528 16820 74592
rect 16884 74528 16900 74592
rect 16964 74528 16980 74592
rect 17044 74528 17060 74592
rect 17124 74528 17140 74592
rect 17204 74528 17220 74592
rect 17284 74528 17322 74592
rect 16702 74512 17322 74528
rect 16702 74448 16740 74512
rect 16804 74448 16820 74512
rect 16884 74448 16900 74512
rect 16964 74448 16980 74512
rect 17044 74448 17060 74512
rect 17124 74448 17140 74512
rect 17204 74448 17220 74512
rect 17284 74448 17322 74512
rect 16702 74432 17322 74448
rect 16702 74368 16740 74432
rect 16804 74368 16820 74432
rect 16884 74368 16900 74432
rect 16964 74368 16980 74432
rect 17044 74368 17060 74432
rect 17124 74368 17140 74432
rect 17204 74368 17220 74432
rect 17284 74368 17322 74432
rect 16702 74352 17322 74368
rect 16702 74288 16740 74352
rect 16804 74288 16820 74352
rect 16884 74288 16900 74352
rect 16964 74288 16980 74352
rect 17044 74288 17060 74352
rect 17124 74288 17140 74352
rect 17204 74288 17220 74352
rect 17284 74288 17322 74352
rect 16702 64592 17322 74288
rect 16702 64528 16740 64592
rect 16804 64528 16820 64592
rect 16884 64528 16900 64592
rect 16964 64528 16980 64592
rect 17044 64528 17060 64592
rect 17124 64528 17140 64592
rect 17204 64528 17220 64592
rect 17284 64528 17322 64592
rect 16702 64512 17322 64528
rect 16702 64448 16740 64512
rect 16804 64448 16820 64512
rect 16884 64448 16900 64512
rect 16964 64448 16980 64512
rect 17044 64448 17060 64512
rect 17124 64448 17140 64512
rect 17204 64448 17220 64512
rect 17284 64448 17322 64512
rect 16702 64432 17322 64448
rect 16702 64368 16740 64432
rect 16804 64368 16820 64432
rect 16884 64368 16900 64432
rect 16964 64368 16980 64432
rect 17044 64368 17060 64432
rect 17124 64368 17140 64432
rect 17204 64368 17220 64432
rect 17284 64368 17322 64432
rect 16702 64352 17322 64368
rect 16702 64288 16740 64352
rect 16804 64288 16820 64352
rect 16884 64288 16900 64352
rect 16964 64288 16980 64352
rect 17044 64288 17060 64352
rect 17124 64288 17140 64352
rect 17204 64288 17220 64352
rect 17284 64288 17322 64352
rect 16702 54592 17322 64288
rect 16702 54528 16740 54592
rect 16804 54528 16820 54592
rect 16884 54528 16900 54592
rect 16964 54528 16980 54592
rect 17044 54528 17060 54592
rect 17124 54528 17140 54592
rect 17204 54528 17220 54592
rect 17284 54528 17322 54592
rect 16702 54512 17322 54528
rect 16702 54448 16740 54512
rect 16804 54448 16820 54512
rect 16884 54448 16900 54512
rect 16964 54448 16980 54512
rect 17044 54448 17060 54512
rect 17124 54448 17140 54512
rect 17204 54448 17220 54512
rect 17284 54448 17322 54512
rect 16702 54432 17322 54448
rect 16702 54368 16740 54432
rect 16804 54368 16820 54432
rect 16884 54368 16900 54432
rect 16964 54368 16980 54432
rect 17044 54368 17060 54432
rect 17124 54368 17140 54432
rect 17204 54368 17220 54432
rect 17284 54368 17322 54432
rect 16702 54352 17322 54368
rect 16702 54288 16740 54352
rect 16804 54288 16820 54352
rect 16884 54288 16900 54352
rect 16964 54288 16980 54352
rect 17044 54288 17060 54352
rect 17124 54288 17140 54352
rect 17204 54288 17220 54352
rect 17284 54288 17322 54352
rect 16702 44592 17322 54288
rect 16702 44528 16740 44592
rect 16804 44528 16820 44592
rect 16884 44528 16900 44592
rect 16964 44528 16980 44592
rect 17044 44528 17060 44592
rect 17124 44528 17140 44592
rect 17204 44528 17220 44592
rect 17284 44528 17322 44592
rect 16702 44512 17322 44528
rect 16702 44448 16740 44512
rect 16804 44448 16820 44512
rect 16884 44448 16900 44512
rect 16964 44448 16980 44512
rect 17044 44448 17060 44512
rect 17124 44448 17140 44512
rect 17204 44448 17220 44512
rect 17284 44448 17322 44512
rect 16702 44432 17322 44448
rect 16702 44368 16740 44432
rect 16804 44368 16820 44432
rect 16884 44368 16900 44432
rect 16964 44368 16980 44432
rect 17044 44368 17060 44432
rect 17124 44368 17140 44432
rect 17204 44368 17220 44432
rect 17284 44368 17322 44432
rect 16702 44352 17322 44368
rect 16702 44288 16740 44352
rect 16804 44288 16820 44352
rect 16884 44288 16900 44352
rect 16964 44288 16980 44352
rect 17044 44288 17060 44352
rect 17124 44288 17140 44352
rect 17204 44288 17220 44352
rect 17284 44288 17322 44352
rect 16702 34592 17322 44288
rect 16702 34528 16740 34592
rect 16804 34528 16820 34592
rect 16884 34528 16900 34592
rect 16964 34528 16980 34592
rect 17044 34528 17060 34592
rect 17124 34528 17140 34592
rect 17204 34528 17220 34592
rect 17284 34528 17322 34592
rect 16702 34512 17322 34528
rect 16702 34448 16740 34512
rect 16804 34448 16820 34512
rect 16884 34448 16900 34512
rect 16964 34448 16980 34512
rect 17044 34448 17060 34512
rect 17124 34448 17140 34512
rect 17204 34448 17220 34512
rect 17284 34448 17322 34512
rect 16702 34432 17322 34448
rect 16702 34368 16740 34432
rect 16804 34368 16820 34432
rect 16884 34368 16900 34432
rect 16964 34368 16980 34432
rect 17044 34368 17060 34432
rect 17124 34368 17140 34432
rect 17204 34368 17220 34432
rect 17284 34368 17322 34432
rect 16702 34352 17322 34368
rect 16702 34288 16740 34352
rect 16804 34288 16820 34352
rect 16884 34288 16900 34352
rect 16964 34288 16980 34352
rect 17044 34288 17060 34352
rect 17124 34288 17140 34352
rect 17204 34288 17220 34352
rect 17284 34288 17322 34352
rect 16702 24592 17322 34288
rect 16702 24528 16740 24592
rect 16804 24528 16820 24592
rect 16884 24528 16900 24592
rect 16964 24528 16980 24592
rect 17044 24528 17060 24592
rect 17124 24528 17140 24592
rect 17204 24528 17220 24592
rect 17284 24528 17322 24592
rect 16702 24512 17322 24528
rect 16702 24448 16740 24512
rect 16804 24448 16820 24512
rect 16884 24448 16900 24512
rect 16964 24448 16980 24512
rect 17044 24448 17060 24512
rect 17124 24448 17140 24512
rect 17204 24448 17220 24512
rect 17284 24448 17322 24512
rect 16702 24432 17322 24448
rect 16702 24368 16740 24432
rect 16804 24368 16820 24432
rect 16884 24368 16900 24432
rect 16964 24368 16980 24432
rect 17044 24368 17060 24432
rect 17124 24368 17140 24432
rect 17204 24368 17220 24432
rect 17284 24368 17322 24432
rect 16702 24352 17322 24368
rect 16702 24288 16740 24352
rect 16804 24288 16820 24352
rect 16884 24288 16900 24352
rect 16964 24288 16980 24352
rect 17044 24288 17060 24352
rect 17124 24288 17140 24352
rect 17204 24288 17220 24352
rect 17284 24288 17322 24352
rect 16702 14592 17322 24288
rect 16702 14528 16740 14592
rect 16804 14528 16820 14592
rect 16884 14528 16900 14592
rect 16964 14528 16980 14592
rect 17044 14528 17060 14592
rect 17124 14528 17140 14592
rect 17204 14528 17220 14592
rect 17284 14528 17322 14592
rect 16702 14512 17322 14528
rect 16702 14448 16740 14512
rect 16804 14448 16820 14512
rect 16884 14448 16900 14512
rect 16964 14448 16980 14512
rect 17044 14448 17060 14512
rect 17124 14448 17140 14512
rect 17204 14448 17220 14512
rect 17284 14448 17322 14512
rect 16702 14432 17322 14448
rect 16702 14368 16740 14432
rect 16804 14368 16820 14432
rect 16884 14368 16900 14432
rect 16964 14368 16980 14432
rect 17044 14368 17060 14432
rect 17124 14368 17140 14432
rect 17204 14368 17220 14432
rect 17284 14368 17322 14432
rect 16702 14352 17322 14368
rect 16702 14288 16740 14352
rect 16804 14288 16820 14352
rect 16884 14288 16900 14352
rect 16964 14288 16980 14352
rect 17044 14288 17060 14352
rect 17124 14288 17140 14352
rect 17204 14288 17220 14352
rect 17284 14288 17322 14352
rect 16702 4592 17322 14288
rect 16702 4528 16740 4592
rect 16804 4528 16820 4592
rect 16884 4528 16900 4592
rect 16964 4528 16980 4592
rect 17044 4528 17060 4592
rect 17124 4528 17140 4592
rect 17204 4528 17220 4592
rect 17284 4528 17322 4592
rect 16702 4512 17322 4528
rect 16702 4448 16740 4512
rect 16804 4448 16820 4512
rect 16884 4448 16900 4512
rect 16964 4448 16980 4512
rect 17044 4448 17060 4512
rect 17124 4448 17140 4512
rect 17204 4448 17220 4512
rect 17284 4448 17322 4512
rect 16702 4432 17322 4448
rect 16702 4368 16740 4432
rect 16804 4368 16820 4432
rect 16884 4368 16900 4432
rect 16964 4368 16980 4432
rect 17044 4368 17060 4432
rect 17124 4368 17140 4432
rect 17204 4368 17220 4432
rect 17284 4368 17322 4432
rect 16702 4352 17322 4368
rect 16702 4288 16740 4352
rect 16804 4288 16820 4352
rect 16884 4288 16900 4352
rect 16964 4288 16980 4352
rect 17044 4288 17060 4352
rect 17124 4288 17140 4352
rect 17204 4288 17220 4352
rect 17284 4288 17322 4352
rect 16702 0 17322 4288
rect 19702 82240 20322 87000
rect 19702 82176 19740 82240
rect 19804 82176 19820 82240
rect 19884 82176 19900 82240
rect 19964 82176 19980 82240
rect 20044 82176 20060 82240
rect 20124 82176 20140 82240
rect 20204 82176 20220 82240
rect 20284 82176 20322 82240
rect 19702 82160 20322 82176
rect 19702 82096 19740 82160
rect 19804 82096 19820 82160
rect 19884 82096 19900 82160
rect 19964 82096 19980 82160
rect 20044 82096 20060 82160
rect 20124 82096 20140 82160
rect 20204 82096 20220 82160
rect 20284 82096 20322 82160
rect 19702 82080 20322 82096
rect 19702 82016 19740 82080
rect 19804 82016 19820 82080
rect 19884 82016 19900 82080
rect 19964 82016 19980 82080
rect 20044 82016 20060 82080
rect 20124 82016 20140 82080
rect 20204 82016 20220 82080
rect 20284 82016 20322 82080
rect 19702 82000 20322 82016
rect 19702 81936 19740 82000
rect 19804 81936 19820 82000
rect 19884 81936 19900 82000
rect 19964 81936 19980 82000
rect 20044 81936 20060 82000
rect 20124 81936 20140 82000
rect 20204 81936 20220 82000
rect 20284 81936 20322 82000
rect 19702 72240 20322 81936
rect 19702 72176 19740 72240
rect 19804 72176 19820 72240
rect 19884 72176 19900 72240
rect 19964 72176 19980 72240
rect 20044 72176 20060 72240
rect 20124 72176 20140 72240
rect 20204 72176 20220 72240
rect 20284 72176 20322 72240
rect 19702 72160 20322 72176
rect 19702 72096 19740 72160
rect 19804 72096 19820 72160
rect 19884 72096 19900 72160
rect 19964 72096 19980 72160
rect 20044 72096 20060 72160
rect 20124 72096 20140 72160
rect 20204 72096 20220 72160
rect 20284 72096 20322 72160
rect 19702 72080 20322 72096
rect 19702 72016 19740 72080
rect 19804 72016 19820 72080
rect 19884 72016 19900 72080
rect 19964 72016 19980 72080
rect 20044 72016 20060 72080
rect 20124 72016 20140 72080
rect 20204 72016 20220 72080
rect 20284 72016 20322 72080
rect 19702 72000 20322 72016
rect 19702 71936 19740 72000
rect 19804 71936 19820 72000
rect 19884 71936 19900 72000
rect 19964 71936 19980 72000
rect 20044 71936 20060 72000
rect 20124 71936 20140 72000
rect 20204 71936 20220 72000
rect 20284 71936 20322 72000
rect 19702 62240 20322 71936
rect 19702 62176 19740 62240
rect 19804 62176 19820 62240
rect 19884 62176 19900 62240
rect 19964 62176 19980 62240
rect 20044 62176 20060 62240
rect 20124 62176 20140 62240
rect 20204 62176 20220 62240
rect 20284 62176 20322 62240
rect 19702 62160 20322 62176
rect 19702 62096 19740 62160
rect 19804 62096 19820 62160
rect 19884 62096 19900 62160
rect 19964 62096 19980 62160
rect 20044 62096 20060 62160
rect 20124 62096 20140 62160
rect 20204 62096 20220 62160
rect 20284 62096 20322 62160
rect 19702 62080 20322 62096
rect 19702 62016 19740 62080
rect 19804 62016 19820 62080
rect 19884 62016 19900 62080
rect 19964 62016 19980 62080
rect 20044 62016 20060 62080
rect 20124 62016 20140 62080
rect 20204 62016 20220 62080
rect 20284 62016 20322 62080
rect 19702 62000 20322 62016
rect 19702 61936 19740 62000
rect 19804 61936 19820 62000
rect 19884 61936 19900 62000
rect 19964 61936 19980 62000
rect 20044 61936 20060 62000
rect 20124 61936 20140 62000
rect 20204 61936 20220 62000
rect 20284 61936 20322 62000
rect 19702 52240 20322 61936
rect 19702 52176 19740 52240
rect 19804 52176 19820 52240
rect 19884 52176 19900 52240
rect 19964 52176 19980 52240
rect 20044 52176 20060 52240
rect 20124 52176 20140 52240
rect 20204 52176 20220 52240
rect 20284 52176 20322 52240
rect 19702 52160 20322 52176
rect 19702 52096 19740 52160
rect 19804 52096 19820 52160
rect 19884 52096 19900 52160
rect 19964 52096 19980 52160
rect 20044 52096 20060 52160
rect 20124 52096 20140 52160
rect 20204 52096 20220 52160
rect 20284 52096 20322 52160
rect 19702 52080 20322 52096
rect 19702 52016 19740 52080
rect 19804 52016 19820 52080
rect 19884 52016 19900 52080
rect 19964 52016 19980 52080
rect 20044 52016 20060 52080
rect 20124 52016 20140 52080
rect 20204 52016 20220 52080
rect 20284 52016 20322 52080
rect 19702 52000 20322 52016
rect 19702 51936 19740 52000
rect 19804 51936 19820 52000
rect 19884 51936 19900 52000
rect 19964 51936 19980 52000
rect 20044 51936 20060 52000
rect 20124 51936 20140 52000
rect 20204 51936 20220 52000
rect 20284 51936 20322 52000
rect 19702 42240 20322 51936
rect 19702 42176 19740 42240
rect 19804 42176 19820 42240
rect 19884 42176 19900 42240
rect 19964 42176 19980 42240
rect 20044 42176 20060 42240
rect 20124 42176 20140 42240
rect 20204 42176 20220 42240
rect 20284 42176 20322 42240
rect 19702 42160 20322 42176
rect 19702 42096 19740 42160
rect 19804 42096 19820 42160
rect 19884 42096 19900 42160
rect 19964 42096 19980 42160
rect 20044 42096 20060 42160
rect 20124 42096 20140 42160
rect 20204 42096 20220 42160
rect 20284 42096 20322 42160
rect 19702 42080 20322 42096
rect 19702 42016 19740 42080
rect 19804 42016 19820 42080
rect 19884 42016 19900 42080
rect 19964 42016 19980 42080
rect 20044 42016 20060 42080
rect 20124 42016 20140 42080
rect 20204 42016 20220 42080
rect 20284 42016 20322 42080
rect 19702 42000 20322 42016
rect 19702 41936 19740 42000
rect 19804 41936 19820 42000
rect 19884 41936 19900 42000
rect 19964 41936 19980 42000
rect 20044 41936 20060 42000
rect 20124 41936 20140 42000
rect 20204 41936 20220 42000
rect 20284 41936 20322 42000
rect 19702 32240 20322 41936
rect 19702 32176 19740 32240
rect 19804 32176 19820 32240
rect 19884 32176 19900 32240
rect 19964 32176 19980 32240
rect 20044 32176 20060 32240
rect 20124 32176 20140 32240
rect 20204 32176 20220 32240
rect 20284 32176 20322 32240
rect 19702 32160 20322 32176
rect 19702 32096 19740 32160
rect 19804 32096 19820 32160
rect 19884 32096 19900 32160
rect 19964 32096 19980 32160
rect 20044 32096 20060 32160
rect 20124 32096 20140 32160
rect 20204 32096 20220 32160
rect 20284 32096 20322 32160
rect 19702 32080 20322 32096
rect 19702 32016 19740 32080
rect 19804 32016 19820 32080
rect 19884 32016 19900 32080
rect 19964 32016 19980 32080
rect 20044 32016 20060 32080
rect 20124 32016 20140 32080
rect 20204 32016 20220 32080
rect 20284 32016 20322 32080
rect 19702 32000 20322 32016
rect 19702 31936 19740 32000
rect 19804 31936 19820 32000
rect 19884 31936 19900 32000
rect 19964 31936 19980 32000
rect 20044 31936 20060 32000
rect 20124 31936 20140 32000
rect 20204 31936 20220 32000
rect 20284 31936 20322 32000
rect 19702 22240 20322 31936
rect 19702 22176 19740 22240
rect 19804 22176 19820 22240
rect 19884 22176 19900 22240
rect 19964 22176 19980 22240
rect 20044 22176 20060 22240
rect 20124 22176 20140 22240
rect 20204 22176 20220 22240
rect 20284 22176 20322 22240
rect 19702 22160 20322 22176
rect 19702 22096 19740 22160
rect 19804 22096 19820 22160
rect 19884 22096 19900 22160
rect 19964 22096 19980 22160
rect 20044 22096 20060 22160
rect 20124 22096 20140 22160
rect 20204 22096 20220 22160
rect 20284 22096 20322 22160
rect 19702 22080 20322 22096
rect 19702 22016 19740 22080
rect 19804 22016 19820 22080
rect 19884 22016 19900 22080
rect 19964 22016 19980 22080
rect 20044 22016 20060 22080
rect 20124 22016 20140 22080
rect 20204 22016 20220 22080
rect 20284 22016 20322 22080
rect 19702 22000 20322 22016
rect 19702 21936 19740 22000
rect 19804 21936 19820 22000
rect 19884 21936 19900 22000
rect 19964 21936 19980 22000
rect 20044 21936 20060 22000
rect 20124 21936 20140 22000
rect 20204 21936 20220 22000
rect 20284 21936 20322 22000
rect 19702 12240 20322 21936
rect 19702 12176 19740 12240
rect 19804 12176 19820 12240
rect 19884 12176 19900 12240
rect 19964 12176 19980 12240
rect 20044 12176 20060 12240
rect 20124 12176 20140 12240
rect 20204 12176 20220 12240
rect 20284 12176 20322 12240
rect 19702 12160 20322 12176
rect 19702 12096 19740 12160
rect 19804 12096 19820 12160
rect 19884 12096 19900 12160
rect 19964 12096 19980 12160
rect 20044 12096 20060 12160
rect 20124 12096 20140 12160
rect 20204 12096 20220 12160
rect 20284 12096 20322 12160
rect 19702 12080 20322 12096
rect 19702 12016 19740 12080
rect 19804 12016 19820 12080
rect 19884 12016 19900 12080
rect 19964 12016 19980 12080
rect 20044 12016 20060 12080
rect 20124 12016 20140 12080
rect 20204 12016 20220 12080
rect 20284 12016 20322 12080
rect 19702 12000 20322 12016
rect 19702 11936 19740 12000
rect 19804 11936 19820 12000
rect 19884 11936 19900 12000
rect 19964 11936 19980 12000
rect 20044 11936 20060 12000
rect 20124 11936 20140 12000
rect 20204 11936 20220 12000
rect 20284 11936 20322 12000
rect 19702 2240 20322 11936
rect 19702 2176 19740 2240
rect 19804 2176 19820 2240
rect 19884 2176 19900 2240
rect 19964 2176 19980 2240
rect 20044 2176 20060 2240
rect 20124 2176 20140 2240
rect 20204 2176 20220 2240
rect 20284 2176 20322 2240
rect 19702 2160 20322 2176
rect 19702 2096 19740 2160
rect 19804 2096 19820 2160
rect 19884 2096 19900 2160
rect 19964 2096 19980 2160
rect 20044 2096 20060 2160
rect 20124 2096 20140 2160
rect 20204 2096 20220 2160
rect 20284 2096 20322 2160
rect 19702 2080 20322 2096
rect 19702 2016 19740 2080
rect 19804 2016 19820 2080
rect 19884 2016 19900 2080
rect 19964 2016 19980 2080
rect 20044 2016 20060 2080
rect 20124 2016 20140 2080
rect 20204 2016 20220 2080
rect 20284 2016 20322 2080
rect 19702 2000 20322 2016
rect 19702 1936 19740 2000
rect 19804 1936 19820 2000
rect 19884 1936 19900 2000
rect 19964 1936 19980 2000
rect 20044 1936 20060 2000
rect 20124 1936 20140 2000
rect 20204 1936 20220 2000
rect 20284 1936 20322 2000
rect 19702 0 20322 1936
rect 22702 84592 23322 87000
rect 22702 84528 22740 84592
rect 22804 84528 22820 84592
rect 22884 84528 22900 84592
rect 22964 84528 22980 84592
rect 23044 84528 23060 84592
rect 23124 84528 23140 84592
rect 23204 84528 23220 84592
rect 23284 84528 23322 84592
rect 22702 84512 23322 84528
rect 22702 84448 22740 84512
rect 22804 84448 22820 84512
rect 22884 84448 22900 84512
rect 22964 84448 22980 84512
rect 23044 84448 23060 84512
rect 23124 84448 23140 84512
rect 23204 84448 23220 84512
rect 23284 84448 23322 84512
rect 22702 84432 23322 84448
rect 22702 84368 22740 84432
rect 22804 84368 22820 84432
rect 22884 84368 22900 84432
rect 22964 84368 22980 84432
rect 23044 84368 23060 84432
rect 23124 84368 23140 84432
rect 23204 84368 23220 84432
rect 23284 84368 23322 84432
rect 22702 84352 23322 84368
rect 22702 84288 22740 84352
rect 22804 84288 22820 84352
rect 22884 84288 22900 84352
rect 22964 84288 22980 84352
rect 23044 84288 23060 84352
rect 23124 84288 23140 84352
rect 23204 84288 23220 84352
rect 23284 84288 23322 84352
rect 22702 74592 23322 84288
rect 22702 74528 22740 74592
rect 22804 74528 22820 74592
rect 22884 74528 22900 74592
rect 22964 74528 22980 74592
rect 23044 74528 23060 74592
rect 23124 74528 23140 74592
rect 23204 74528 23220 74592
rect 23284 74528 23322 74592
rect 22702 74512 23322 74528
rect 22702 74448 22740 74512
rect 22804 74448 22820 74512
rect 22884 74448 22900 74512
rect 22964 74448 22980 74512
rect 23044 74448 23060 74512
rect 23124 74448 23140 74512
rect 23204 74448 23220 74512
rect 23284 74448 23322 74512
rect 22702 74432 23322 74448
rect 22702 74368 22740 74432
rect 22804 74368 22820 74432
rect 22884 74368 22900 74432
rect 22964 74368 22980 74432
rect 23044 74368 23060 74432
rect 23124 74368 23140 74432
rect 23204 74368 23220 74432
rect 23284 74368 23322 74432
rect 22702 74352 23322 74368
rect 22702 74288 22740 74352
rect 22804 74288 22820 74352
rect 22884 74288 22900 74352
rect 22964 74288 22980 74352
rect 23044 74288 23060 74352
rect 23124 74288 23140 74352
rect 23204 74288 23220 74352
rect 23284 74288 23322 74352
rect 22702 64592 23322 74288
rect 22702 64528 22740 64592
rect 22804 64528 22820 64592
rect 22884 64528 22900 64592
rect 22964 64528 22980 64592
rect 23044 64528 23060 64592
rect 23124 64528 23140 64592
rect 23204 64528 23220 64592
rect 23284 64528 23322 64592
rect 22702 64512 23322 64528
rect 22702 64448 22740 64512
rect 22804 64448 22820 64512
rect 22884 64448 22900 64512
rect 22964 64448 22980 64512
rect 23044 64448 23060 64512
rect 23124 64448 23140 64512
rect 23204 64448 23220 64512
rect 23284 64448 23322 64512
rect 22702 64432 23322 64448
rect 22702 64368 22740 64432
rect 22804 64368 22820 64432
rect 22884 64368 22900 64432
rect 22964 64368 22980 64432
rect 23044 64368 23060 64432
rect 23124 64368 23140 64432
rect 23204 64368 23220 64432
rect 23284 64368 23322 64432
rect 22702 64352 23322 64368
rect 22702 64288 22740 64352
rect 22804 64288 22820 64352
rect 22884 64288 22900 64352
rect 22964 64288 22980 64352
rect 23044 64288 23060 64352
rect 23124 64288 23140 64352
rect 23204 64288 23220 64352
rect 23284 64288 23322 64352
rect 22702 54592 23322 64288
rect 22702 54528 22740 54592
rect 22804 54528 22820 54592
rect 22884 54528 22900 54592
rect 22964 54528 22980 54592
rect 23044 54528 23060 54592
rect 23124 54528 23140 54592
rect 23204 54528 23220 54592
rect 23284 54528 23322 54592
rect 22702 54512 23322 54528
rect 22702 54448 22740 54512
rect 22804 54448 22820 54512
rect 22884 54448 22900 54512
rect 22964 54448 22980 54512
rect 23044 54448 23060 54512
rect 23124 54448 23140 54512
rect 23204 54448 23220 54512
rect 23284 54448 23322 54512
rect 22702 54432 23322 54448
rect 22702 54368 22740 54432
rect 22804 54368 22820 54432
rect 22884 54368 22900 54432
rect 22964 54368 22980 54432
rect 23044 54368 23060 54432
rect 23124 54368 23140 54432
rect 23204 54368 23220 54432
rect 23284 54368 23322 54432
rect 22702 54352 23322 54368
rect 22702 54288 22740 54352
rect 22804 54288 22820 54352
rect 22884 54288 22900 54352
rect 22964 54288 22980 54352
rect 23044 54288 23060 54352
rect 23124 54288 23140 54352
rect 23204 54288 23220 54352
rect 23284 54288 23322 54352
rect 22702 44592 23322 54288
rect 22702 44528 22740 44592
rect 22804 44528 22820 44592
rect 22884 44528 22900 44592
rect 22964 44528 22980 44592
rect 23044 44528 23060 44592
rect 23124 44528 23140 44592
rect 23204 44528 23220 44592
rect 23284 44528 23322 44592
rect 22702 44512 23322 44528
rect 22702 44448 22740 44512
rect 22804 44448 22820 44512
rect 22884 44448 22900 44512
rect 22964 44448 22980 44512
rect 23044 44448 23060 44512
rect 23124 44448 23140 44512
rect 23204 44448 23220 44512
rect 23284 44448 23322 44512
rect 22702 44432 23322 44448
rect 22702 44368 22740 44432
rect 22804 44368 22820 44432
rect 22884 44368 22900 44432
rect 22964 44368 22980 44432
rect 23044 44368 23060 44432
rect 23124 44368 23140 44432
rect 23204 44368 23220 44432
rect 23284 44368 23322 44432
rect 22702 44352 23322 44368
rect 22702 44288 22740 44352
rect 22804 44288 22820 44352
rect 22884 44288 22900 44352
rect 22964 44288 22980 44352
rect 23044 44288 23060 44352
rect 23124 44288 23140 44352
rect 23204 44288 23220 44352
rect 23284 44288 23322 44352
rect 22702 34592 23322 44288
rect 22702 34528 22740 34592
rect 22804 34528 22820 34592
rect 22884 34528 22900 34592
rect 22964 34528 22980 34592
rect 23044 34528 23060 34592
rect 23124 34528 23140 34592
rect 23204 34528 23220 34592
rect 23284 34528 23322 34592
rect 22702 34512 23322 34528
rect 22702 34448 22740 34512
rect 22804 34448 22820 34512
rect 22884 34448 22900 34512
rect 22964 34448 22980 34512
rect 23044 34448 23060 34512
rect 23124 34448 23140 34512
rect 23204 34448 23220 34512
rect 23284 34448 23322 34512
rect 22702 34432 23322 34448
rect 22702 34368 22740 34432
rect 22804 34368 22820 34432
rect 22884 34368 22900 34432
rect 22964 34368 22980 34432
rect 23044 34368 23060 34432
rect 23124 34368 23140 34432
rect 23204 34368 23220 34432
rect 23284 34368 23322 34432
rect 22702 34352 23322 34368
rect 22702 34288 22740 34352
rect 22804 34288 22820 34352
rect 22884 34288 22900 34352
rect 22964 34288 22980 34352
rect 23044 34288 23060 34352
rect 23124 34288 23140 34352
rect 23204 34288 23220 34352
rect 23284 34288 23322 34352
rect 22702 24592 23322 34288
rect 22702 24528 22740 24592
rect 22804 24528 22820 24592
rect 22884 24528 22900 24592
rect 22964 24528 22980 24592
rect 23044 24528 23060 24592
rect 23124 24528 23140 24592
rect 23204 24528 23220 24592
rect 23284 24528 23322 24592
rect 22702 24512 23322 24528
rect 22702 24448 22740 24512
rect 22804 24448 22820 24512
rect 22884 24448 22900 24512
rect 22964 24448 22980 24512
rect 23044 24448 23060 24512
rect 23124 24448 23140 24512
rect 23204 24448 23220 24512
rect 23284 24448 23322 24512
rect 22702 24432 23322 24448
rect 22702 24368 22740 24432
rect 22804 24368 22820 24432
rect 22884 24368 22900 24432
rect 22964 24368 22980 24432
rect 23044 24368 23060 24432
rect 23124 24368 23140 24432
rect 23204 24368 23220 24432
rect 23284 24368 23322 24432
rect 22702 24352 23322 24368
rect 22702 24288 22740 24352
rect 22804 24288 22820 24352
rect 22884 24288 22900 24352
rect 22964 24288 22980 24352
rect 23044 24288 23060 24352
rect 23124 24288 23140 24352
rect 23204 24288 23220 24352
rect 23284 24288 23322 24352
rect 22702 14592 23322 24288
rect 22702 14528 22740 14592
rect 22804 14528 22820 14592
rect 22884 14528 22900 14592
rect 22964 14528 22980 14592
rect 23044 14528 23060 14592
rect 23124 14528 23140 14592
rect 23204 14528 23220 14592
rect 23284 14528 23322 14592
rect 22702 14512 23322 14528
rect 22702 14448 22740 14512
rect 22804 14448 22820 14512
rect 22884 14448 22900 14512
rect 22964 14448 22980 14512
rect 23044 14448 23060 14512
rect 23124 14448 23140 14512
rect 23204 14448 23220 14512
rect 23284 14448 23322 14512
rect 22702 14432 23322 14448
rect 22702 14368 22740 14432
rect 22804 14368 22820 14432
rect 22884 14368 22900 14432
rect 22964 14368 22980 14432
rect 23044 14368 23060 14432
rect 23124 14368 23140 14432
rect 23204 14368 23220 14432
rect 23284 14368 23322 14432
rect 22702 14352 23322 14368
rect 22702 14288 22740 14352
rect 22804 14288 22820 14352
rect 22884 14288 22900 14352
rect 22964 14288 22980 14352
rect 23044 14288 23060 14352
rect 23124 14288 23140 14352
rect 23204 14288 23220 14352
rect 23284 14288 23322 14352
rect 22702 4592 23322 14288
rect 22702 4528 22740 4592
rect 22804 4528 22820 4592
rect 22884 4528 22900 4592
rect 22964 4528 22980 4592
rect 23044 4528 23060 4592
rect 23124 4528 23140 4592
rect 23204 4528 23220 4592
rect 23284 4528 23322 4592
rect 22702 4512 23322 4528
rect 22702 4448 22740 4512
rect 22804 4448 22820 4512
rect 22884 4448 22900 4512
rect 22964 4448 22980 4512
rect 23044 4448 23060 4512
rect 23124 4448 23140 4512
rect 23204 4448 23220 4512
rect 23284 4448 23322 4512
rect 22702 4432 23322 4448
rect 22702 4368 22740 4432
rect 22804 4368 22820 4432
rect 22884 4368 22900 4432
rect 22964 4368 22980 4432
rect 23044 4368 23060 4432
rect 23124 4368 23140 4432
rect 23204 4368 23220 4432
rect 23284 4368 23322 4432
rect 22702 4352 23322 4368
rect 22702 4288 22740 4352
rect 22804 4288 22820 4352
rect 22884 4288 22900 4352
rect 22964 4288 22980 4352
rect 23044 4288 23060 4352
rect 23124 4288 23140 4352
rect 23204 4288 23220 4352
rect 23284 4288 23322 4352
rect 22702 0 23322 4288
rect 25702 82240 26322 87000
rect 25702 82176 25740 82240
rect 25804 82176 25820 82240
rect 25884 82176 25900 82240
rect 25964 82176 25980 82240
rect 26044 82176 26060 82240
rect 26124 82176 26140 82240
rect 26204 82176 26220 82240
rect 26284 82176 26322 82240
rect 25702 82160 26322 82176
rect 25702 82096 25740 82160
rect 25804 82096 25820 82160
rect 25884 82096 25900 82160
rect 25964 82096 25980 82160
rect 26044 82096 26060 82160
rect 26124 82096 26140 82160
rect 26204 82096 26220 82160
rect 26284 82096 26322 82160
rect 25702 82080 26322 82096
rect 25702 82016 25740 82080
rect 25804 82016 25820 82080
rect 25884 82016 25900 82080
rect 25964 82016 25980 82080
rect 26044 82016 26060 82080
rect 26124 82016 26140 82080
rect 26204 82016 26220 82080
rect 26284 82016 26322 82080
rect 25702 82000 26322 82016
rect 25702 81936 25740 82000
rect 25804 81936 25820 82000
rect 25884 81936 25900 82000
rect 25964 81936 25980 82000
rect 26044 81936 26060 82000
rect 26124 81936 26140 82000
rect 26204 81936 26220 82000
rect 26284 81936 26322 82000
rect 25702 72240 26322 81936
rect 25702 72176 25740 72240
rect 25804 72176 25820 72240
rect 25884 72176 25900 72240
rect 25964 72176 25980 72240
rect 26044 72176 26060 72240
rect 26124 72176 26140 72240
rect 26204 72176 26220 72240
rect 26284 72176 26322 72240
rect 25702 72160 26322 72176
rect 25702 72096 25740 72160
rect 25804 72096 25820 72160
rect 25884 72096 25900 72160
rect 25964 72096 25980 72160
rect 26044 72096 26060 72160
rect 26124 72096 26140 72160
rect 26204 72096 26220 72160
rect 26284 72096 26322 72160
rect 25702 72080 26322 72096
rect 25702 72016 25740 72080
rect 25804 72016 25820 72080
rect 25884 72016 25900 72080
rect 25964 72016 25980 72080
rect 26044 72016 26060 72080
rect 26124 72016 26140 72080
rect 26204 72016 26220 72080
rect 26284 72016 26322 72080
rect 25702 72000 26322 72016
rect 25702 71936 25740 72000
rect 25804 71936 25820 72000
rect 25884 71936 25900 72000
rect 25964 71936 25980 72000
rect 26044 71936 26060 72000
rect 26124 71936 26140 72000
rect 26204 71936 26220 72000
rect 26284 71936 26322 72000
rect 25702 62240 26322 71936
rect 25702 62176 25740 62240
rect 25804 62176 25820 62240
rect 25884 62176 25900 62240
rect 25964 62176 25980 62240
rect 26044 62176 26060 62240
rect 26124 62176 26140 62240
rect 26204 62176 26220 62240
rect 26284 62176 26322 62240
rect 25702 62160 26322 62176
rect 25702 62096 25740 62160
rect 25804 62096 25820 62160
rect 25884 62096 25900 62160
rect 25964 62096 25980 62160
rect 26044 62096 26060 62160
rect 26124 62096 26140 62160
rect 26204 62096 26220 62160
rect 26284 62096 26322 62160
rect 25702 62080 26322 62096
rect 25702 62016 25740 62080
rect 25804 62016 25820 62080
rect 25884 62016 25900 62080
rect 25964 62016 25980 62080
rect 26044 62016 26060 62080
rect 26124 62016 26140 62080
rect 26204 62016 26220 62080
rect 26284 62016 26322 62080
rect 25702 62000 26322 62016
rect 25702 61936 25740 62000
rect 25804 61936 25820 62000
rect 25884 61936 25900 62000
rect 25964 61936 25980 62000
rect 26044 61936 26060 62000
rect 26124 61936 26140 62000
rect 26204 61936 26220 62000
rect 26284 61936 26322 62000
rect 25702 52240 26322 61936
rect 25702 52176 25740 52240
rect 25804 52176 25820 52240
rect 25884 52176 25900 52240
rect 25964 52176 25980 52240
rect 26044 52176 26060 52240
rect 26124 52176 26140 52240
rect 26204 52176 26220 52240
rect 26284 52176 26322 52240
rect 25702 52160 26322 52176
rect 25702 52096 25740 52160
rect 25804 52096 25820 52160
rect 25884 52096 25900 52160
rect 25964 52096 25980 52160
rect 26044 52096 26060 52160
rect 26124 52096 26140 52160
rect 26204 52096 26220 52160
rect 26284 52096 26322 52160
rect 25702 52080 26322 52096
rect 25702 52016 25740 52080
rect 25804 52016 25820 52080
rect 25884 52016 25900 52080
rect 25964 52016 25980 52080
rect 26044 52016 26060 52080
rect 26124 52016 26140 52080
rect 26204 52016 26220 52080
rect 26284 52016 26322 52080
rect 25702 52000 26322 52016
rect 25702 51936 25740 52000
rect 25804 51936 25820 52000
rect 25884 51936 25900 52000
rect 25964 51936 25980 52000
rect 26044 51936 26060 52000
rect 26124 51936 26140 52000
rect 26204 51936 26220 52000
rect 26284 51936 26322 52000
rect 25702 42240 26322 51936
rect 25702 42176 25740 42240
rect 25804 42176 25820 42240
rect 25884 42176 25900 42240
rect 25964 42176 25980 42240
rect 26044 42176 26060 42240
rect 26124 42176 26140 42240
rect 26204 42176 26220 42240
rect 26284 42176 26322 42240
rect 25702 42160 26322 42176
rect 25702 42096 25740 42160
rect 25804 42096 25820 42160
rect 25884 42096 25900 42160
rect 25964 42096 25980 42160
rect 26044 42096 26060 42160
rect 26124 42096 26140 42160
rect 26204 42096 26220 42160
rect 26284 42096 26322 42160
rect 25702 42080 26322 42096
rect 25702 42016 25740 42080
rect 25804 42016 25820 42080
rect 25884 42016 25900 42080
rect 25964 42016 25980 42080
rect 26044 42016 26060 42080
rect 26124 42016 26140 42080
rect 26204 42016 26220 42080
rect 26284 42016 26322 42080
rect 25702 42000 26322 42016
rect 25702 41936 25740 42000
rect 25804 41936 25820 42000
rect 25884 41936 25900 42000
rect 25964 41936 25980 42000
rect 26044 41936 26060 42000
rect 26124 41936 26140 42000
rect 26204 41936 26220 42000
rect 26284 41936 26322 42000
rect 25702 32240 26322 41936
rect 25702 32176 25740 32240
rect 25804 32176 25820 32240
rect 25884 32176 25900 32240
rect 25964 32176 25980 32240
rect 26044 32176 26060 32240
rect 26124 32176 26140 32240
rect 26204 32176 26220 32240
rect 26284 32176 26322 32240
rect 25702 32160 26322 32176
rect 25702 32096 25740 32160
rect 25804 32096 25820 32160
rect 25884 32096 25900 32160
rect 25964 32096 25980 32160
rect 26044 32096 26060 32160
rect 26124 32096 26140 32160
rect 26204 32096 26220 32160
rect 26284 32096 26322 32160
rect 25702 32080 26322 32096
rect 25702 32016 25740 32080
rect 25804 32016 25820 32080
rect 25884 32016 25900 32080
rect 25964 32016 25980 32080
rect 26044 32016 26060 32080
rect 26124 32016 26140 32080
rect 26204 32016 26220 32080
rect 26284 32016 26322 32080
rect 25702 32000 26322 32016
rect 25702 31936 25740 32000
rect 25804 31936 25820 32000
rect 25884 31936 25900 32000
rect 25964 31936 25980 32000
rect 26044 31936 26060 32000
rect 26124 31936 26140 32000
rect 26204 31936 26220 32000
rect 26284 31936 26322 32000
rect 25702 22240 26322 31936
rect 25702 22176 25740 22240
rect 25804 22176 25820 22240
rect 25884 22176 25900 22240
rect 25964 22176 25980 22240
rect 26044 22176 26060 22240
rect 26124 22176 26140 22240
rect 26204 22176 26220 22240
rect 26284 22176 26322 22240
rect 25702 22160 26322 22176
rect 25702 22096 25740 22160
rect 25804 22096 25820 22160
rect 25884 22096 25900 22160
rect 25964 22096 25980 22160
rect 26044 22096 26060 22160
rect 26124 22096 26140 22160
rect 26204 22096 26220 22160
rect 26284 22096 26322 22160
rect 25702 22080 26322 22096
rect 25702 22016 25740 22080
rect 25804 22016 25820 22080
rect 25884 22016 25900 22080
rect 25964 22016 25980 22080
rect 26044 22016 26060 22080
rect 26124 22016 26140 22080
rect 26204 22016 26220 22080
rect 26284 22016 26322 22080
rect 25702 22000 26322 22016
rect 25702 21936 25740 22000
rect 25804 21936 25820 22000
rect 25884 21936 25900 22000
rect 25964 21936 25980 22000
rect 26044 21936 26060 22000
rect 26124 21936 26140 22000
rect 26204 21936 26220 22000
rect 26284 21936 26322 22000
rect 25702 12240 26322 21936
rect 25702 12176 25740 12240
rect 25804 12176 25820 12240
rect 25884 12176 25900 12240
rect 25964 12176 25980 12240
rect 26044 12176 26060 12240
rect 26124 12176 26140 12240
rect 26204 12176 26220 12240
rect 26284 12176 26322 12240
rect 25702 12160 26322 12176
rect 25702 12096 25740 12160
rect 25804 12096 25820 12160
rect 25884 12096 25900 12160
rect 25964 12096 25980 12160
rect 26044 12096 26060 12160
rect 26124 12096 26140 12160
rect 26204 12096 26220 12160
rect 26284 12096 26322 12160
rect 25702 12080 26322 12096
rect 25702 12016 25740 12080
rect 25804 12016 25820 12080
rect 25884 12016 25900 12080
rect 25964 12016 25980 12080
rect 26044 12016 26060 12080
rect 26124 12016 26140 12080
rect 26204 12016 26220 12080
rect 26284 12016 26322 12080
rect 25702 12000 26322 12016
rect 25702 11936 25740 12000
rect 25804 11936 25820 12000
rect 25884 11936 25900 12000
rect 25964 11936 25980 12000
rect 26044 11936 26060 12000
rect 26124 11936 26140 12000
rect 26204 11936 26220 12000
rect 26284 11936 26322 12000
rect 25702 2240 26322 11936
rect 25702 2176 25740 2240
rect 25804 2176 25820 2240
rect 25884 2176 25900 2240
rect 25964 2176 25980 2240
rect 26044 2176 26060 2240
rect 26124 2176 26140 2240
rect 26204 2176 26220 2240
rect 26284 2176 26322 2240
rect 25702 2160 26322 2176
rect 25702 2096 25740 2160
rect 25804 2096 25820 2160
rect 25884 2096 25900 2160
rect 25964 2096 25980 2160
rect 26044 2096 26060 2160
rect 26124 2096 26140 2160
rect 26204 2096 26220 2160
rect 26284 2096 26322 2160
rect 25702 2080 26322 2096
rect 25702 2016 25740 2080
rect 25804 2016 25820 2080
rect 25884 2016 25900 2080
rect 25964 2016 25980 2080
rect 26044 2016 26060 2080
rect 26124 2016 26140 2080
rect 26204 2016 26220 2080
rect 26284 2016 26322 2080
rect 25702 2000 26322 2016
rect 25702 1936 25740 2000
rect 25804 1936 25820 2000
rect 25884 1936 25900 2000
rect 25964 1936 25980 2000
rect 26044 1936 26060 2000
rect 26124 1936 26140 2000
rect 26204 1936 26220 2000
rect 26284 1936 26322 2000
rect 25702 0 26322 1936
rect 28702 84592 29322 87000
rect 28702 84528 28740 84592
rect 28804 84528 28820 84592
rect 28884 84528 28900 84592
rect 28964 84528 28980 84592
rect 29044 84528 29060 84592
rect 29124 84528 29140 84592
rect 29204 84528 29220 84592
rect 29284 84528 29322 84592
rect 28702 84512 29322 84528
rect 28702 84448 28740 84512
rect 28804 84448 28820 84512
rect 28884 84448 28900 84512
rect 28964 84448 28980 84512
rect 29044 84448 29060 84512
rect 29124 84448 29140 84512
rect 29204 84448 29220 84512
rect 29284 84448 29322 84512
rect 28702 84432 29322 84448
rect 28702 84368 28740 84432
rect 28804 84368 28820 84432
rect 28884 84368 28900 84432
rect 28964 84368 28980 84432
rect 29044 84368 29060 84432
rect 29124 84368 29140 84432
rect 29204 84368 29220 84432
rect 29284 84368 29322 84432
rect 28702 84352 29322 84368
rect 28702 84288 28740 84352
rect 28804 84288 28820 84352
rect 28884 84288 28900 84352
rect 28964 84288 28980 84352
rect 29044 84288 29060 84352
rect 29124 84288 29140 84352
rect 29204 84288 29220 84352
rect 29284 84288 29322 84352
rect 28702 74592 29322 84288
rect 28702 74528 28740 74592
rect 28804 74528 28820 74592
rect 28884 74528 28900 74592
rect 28964 74528 28980 74592
rect 29044 74528 29060 74592
rect 29124 74528 29140 74592
rect 29204 74528 29220 74592
rect 29284 74528 29322 74592
rect 28702 74512 29322 74528
rect 28702 74448 28740 74512
rect 28804 74448 28820 74512
rect 28884 74448 28900 74512
rect 28964 74448 28980 74512
rect 29044 74448 29060 74512
rect 29124 74448 29140 74512
rect 29204 74448 29220 74512
rect 29284 74448 29322 74512
rect 28702 74432 29322 74448
rect 28702 74368 28740 74432
rect 28804 74368 28820 74432
rect 28884 74368 28900 74432
rect 28964 74368 28980 74432
rect 29044 74368 29060 74432
rect 29124 74368 29140 74432
rect 29204 74368 29220 74432
rect 29284 74368 29322 74432
rect 28702 74352 29322 74368
rect 28702 74288 28740 74352
rect 28804 74288 28820 74352
rect 28884 74288 28900 74352
rect 28964 74288 28980 74352
rect 29044 74288 29060 74352
rect 29124 74288 29140 74352
rect 29204 74288 29220 74352
rect 29284 74288 29322 74352
rect 28702 64592 29322 74288
rect 28702 64528 28740 64592
rect 28804 64528 28820 64592
rect 28884 64528 28900 64592
rect 28964 64528 28980 64592
rect 29044 64528 29060 64592
rect 29124 64528 29140 64592
rect 29204 64528 29220 64592
rect 29284 64528 29322 64592
rect 28702 64512 29322 64528
rect 28702 64448 28740 64512
rect 28804 64448 28820 64512
rect 28884 64448 28900 64512
rect 28964 64448 28980 64512
rect 29044 64448 29060 64512
rect 29124 64448 29140 64512
rect 29204 64448 29220 64512
rect 29284 64448 29322 64512
rect 28702 64432 29322 64448
rect 28702 64368 28740 64432
rect 28804 64368 28820 64432
rect 28884 64368 28900 64432
rect 28964 64368 28980 64432
rect 29044 64368 29060 64432
rect 29124 64368 29140 64432
rect 29204 64368 29220 64432
rect 29284 64368 29322 64432
rect 28702 64352 29322 64368
rect 28702 64288 28740 64352
rect 28804 64288 28820 64352
rect 28884 64288 28900 64352
rect 28964 64288 28980 64352
rect 29044 64288 29060 64352
rect 29124 64288 29140 64352
rect 29204 64288 29220 64352
rect 29284 64288 29322 64352
rect 28702 54592 29322 64288
rect 28702 54528 28740 54592
rect 28804 54528 28820 54592
rect 28884 54528 28900 54592
rect 28964 54528 28980 54592
rect 29044 54528 29060 54592
rect 29124 54528 29140 54592
rect 29204 54528 29220 54592
rect 29284 54528 29322 54592
rect 28702 54512 29322 54528
rect 28702 54448 28740 54512
rect 28804 54448 28820 54512
rect 28884 54448 28900 54512
rect 28964 54448 28980 54512
rect 29044 54448 29060 54512
rect 29124 54448 29140 54512
rect 29204 54448 29220 54512
rect 29284 54448 29322 54512
rect 28702 54432 29322 54448
rect 28702 54368 28740 54432
rect 28804 54368 28820 54432
rect 28884 54368 28900 54432
rect 28964 54368 28980 54432
rect 29044 54368 29060 54432
rect 29124 54368 29140 54432
rect 29204 54368 29220 54432
rect 29284 54368 29322 54432
rect 28702 54352 29322 54368
rect 28702 54288 28740 54352
rect 28804 54288 28820 54352
rect 28884 54288 28900 54352
rect 28964 54288 28980 54352
rect 29044 54288 29060 54352
rect 29124 54288 29140 54352
rect 29204 54288 29220 54352
rect 29284 54288 29322 54352
rect 28702 44592 29322 54288
rect 28702 44528 28740 44592
rect 28804 44528 28820 44592
rect 28884 44528 28900 44592
rect 28964 44528 28980 44592
rect 29044 44528 29060 44592
rect 29124 44528 29140 44592
rect 29204 44528 29220 44592
rect 29284 44528 29322 44592
rect 28702 44512 29322 44528
rect 28702 44448 28740 44512
rect 28804 44448 28820 44512
rect 28884 44448 28900 44512
rect 28964 44448 28980 44512
rect 29044 44448 29060 44512
rect 29124 44448 29140 44512
rect 29204 44448 29220 44512
rect 29284 44448 29322 44512
rect 28702 44432 29322 44448
rect 28702 44368 28740 44432
rect 28804 44368 28820 44432
rect 28884 44368 28900 44432
rect 28964 44368 28980 44432
rect 29044 44368 29060 44432
rect 29124 44368 29140 44432
rect 29204 44368 29220 44432
rect 29284 44368 29322 44432
rect 28702 44352 29322 44368
rect 28702 44288 28740 44352
rect 28804 44288 28820 44352
rect 28884 44288 28900 44352
rect 28964 44288 28980 44352
rect 29044 44288 29060 44352
rect 29124 44288 29140 44352
rect 29204 44288 29220 44352
rect 29284 44288 29322 44352
rect 28702 34592 29322 44288
rect 28702 34528 28740 34592
rect 28804 34528 28820 34592
rect 28884 34528 28900 34592
rect 28964 34528 28980 34592
rect 29044 34528 29060 34592
rect 29124 34528 29140 34592
rect 29204 34528 29220 34592
rect 29284 34528 29322 34592
rect 28702 34512 29322 34528
rect 28702 34448 28740 34512
rect 28804 34448 28820 34512
rect 28884 34448 28900 34512
rect 28964 34448 28980 34512
rect 29044 34448 29060 34512
rect 29124 34448 29140 34512
rect 29204 34448 29220 34512
rect 29284 34448 29322 34512
rect 28702 34432 29322 34448
rect 28702 34368 28740 34432
rect 28804 34368 28820 34432
rect 28884 34368 28900 34432
rect 28964 34368 28980 34432
rect 29044 34368 29060 34432
rect 29124 34368 29140 34432
rect 29204 34368 29220 34432
rect 29284 34368 29322 34432
rect 28702 34352 29322 34368
rect 28702 34288 28740 34352
rect 28804 34288 28820 34352
rect 28884 34288 28900 34352
rect 28964 34288 28980 34352
rect 29044 34288 29060 34352
rect 29124 34288 29140 34352
rect 29204 34288 29220 34352
rect 29284 34288 29322 34352
rect 28702 24592 29322 34288
rect 28702 24528 28740 24592
rect 28804 24528 28820 24592
rect 28884 24528 28900 24592
rect 28964 24528 28980 24592
rect 29044 24528 29060 24592
rect 29124 24528 29140 24592
rect 29204 24528 29220 24592
rect 29284 24528 29322 24592
rect 28702 24512 29322 24528
rect 28702 24448 28740 24512
rect 28804 24448 28820 24512
rect 28884 24448 28900 24512
rect 28964 24448 28980 24512
rect 29044 24448 29060 24512
rect 29124 24448 29140 24512
rect 29204 24448 29220 24512
rect 29284 24448 29322 24512
rect 28702 24432 29322 24448
rect 28702 24368 28740 24432
rect 28804 24368 28820 24432
rect 28884 24368 28900 24432
rect 28964 24368 28980 24432
rect 29044 24368 29060 24432
rect 29124 24368 29140 24432
rect 29204 24368 29220 24432
rect 29284 24368 29322 24432
rect 28702 24352 29322 24368
rect 28702 24288 28740 24352
rect 28804 24288 28820 24352
rect 28884 24288 28900 24352
rect 28964 24288 28980 24352
rect 29044 24288 29060 24352
rect 29124 24288 29140 24352
rect 29204 24288 29220 24352
rect 29284 24288 29322 24352
rect 28702 14592 29322 24288
rect 28702 14528 28740 14592
rect 28804 14528 28820 14592
rect 28884 14528 28900 14592
rect 28964 14528 28980 14592
rect 29044 14528 29060 14592
rect 29124 14528 29140 14592
rect 29204 14528 29220 14592
rect 29284 14528 29322 14592
rect 28702 14512 29322 14528
rect 28702 14448 28740 14512
rect 28804 14448 28820 14512
rect 28884 14448 28900 14512
rect 28964 14448 28980 14512
rect 29044 14448 29060 14512
rect 29124 14448 29140 14512
rect 29204 14448 29220 14512
rect 29284 14448 29322 14512
rect 28702 14432 29322 14448
rect 28702 14368 28740 14432
rect 28804 14368 28820 14432
rect 28884 14368 28900 14432
rect 28964 14368 28980 14432
rect 29044 14368 29060 14432
rect 29124 14368 29140 14432
rect 29204 14368 29220 14432
rect 29284 14368 29322 14432
rect 28702 14352 29322 14368
rect 28702 14288 28740 14352
rect 28804 14288 28820 14352
rect 28884 14288 28900 14352
rect 28964 14288 28980 14352
rect 29044 14288 29060 14352
rect 29124 14288 29140 14352
rect 29204 14288 29220 14352
rect 29284 14288 29322 14352
rect 28702 4592 29322 14288
rect 28702 4528 28740 4592
rect 28804 4528 28820 4592
rect 28884 4528 28900 4592
rect 28964 4528 28980 4592
rect 29044 4528 29060 4592
rect 29124 4528 29140 4592
rect 29204 4528 29220 4592
rect 29284 4528 29322 4592
rect 28702 4512 29322 4528
rect 28702 4448 28740 4512
rect 28804 4448 28820 4512
rect 28884 4448 28900 4512
rect 28964 4448 28980 4512
rect 29044 4448 29060 4512
rect 29124 4448 29140 4512
rect 29204 4448 29220 4512
rect 29284 4448 29322 4512
rect 28702 4432 29322 4448
rect 28702 4368 28740 4432
rect 28804 4368 28820 4432
rect 28884 4368 28900 4432
rect 28964 4368 28980 4432
rect 29044 4368 29060 4432
rect 29124 4368 29140 4432
rect 29204 4368 29220 4432
rect 29284 4368 29322 4432
rect 28702 4352 29322 4368
rect 28702 4288 28740 4352
rect 28804 4288 28820 4352
rect 28884 4288 28900 4352
rect 28964 4288 28980 4352
rect 29044 4288 29060 4352
rect 29124 4288 29140 4352
rect 29204 4288 29220 4352
rect 29284 4288 29322 4352
rect 28702 0 29322 4288
rect 31702 82240 32322 87000
rect 31702 82176 31740 82240
rect 31804 82176 31820 82240
rect 31884 82176 31900 82240
rect 31964 82176 31980 82240
rect 32044 82176 32060 82240
rect 32124 82176 32140 82240
rect 32204 82176 32220 82240
rect 32284 82176 32322 82240
rect 31702 82160 32322 82176
rect 31702 82096 31740 82160
rect 31804 82096 31820 82160
rect 31884 82096 31900 82160
rect 31964 82096 31980 82160
rect 32044 82096 32060 82160
rect 32124 82096 32140 82160
rect 32204 82096 32220 82160
rect 32284 82096 32322 82160
rect 31702 82080 32322 82096
rect 31702 82016 31740 82080
rect 31804 82016 31820 82080
rect 31884 82016 31900 82080
rect 31964 82016 31980 82080
rect 32044 82016 32060 82080
rect 32124 82016 32140 82080
rect 32204 82016 32220 82080
rect 32284 82016 32322 82080
rect 31702 82000 32322 82016
rect 31702 81936 31740 82000
rect 31804 81936 31820 82000
rect 31884 81936 31900 82000
rect 31964 81936 31980 82000
rect 32044 81936 32060 82000
rect 32124 81936 32140 82000
rect 32204 81936 32220 82000
rect 32284 81936 32322 82000
rect 31702 72240 32322 81936
rect 31702 72176 31740 72240
rect 31804 72176 31820 72240
rect 31884 72176 31900 72240
rect 31964 72176 31980 72240
rect 32044 72176 32060 72240
rect 32124 72176 32140 72240
rect 32204 72176 32220 72240
rect 32284 72176 32322 72240
rect 31702 72160 32322 72176
rect 31702 72096 31740 72160
rect 31804 72096 31820 72160
rect 31884 72096 31900 72160
rect 31964 72096 31980 72160
rect 32044 72096 32060 72160
rect 32124 72096 32140 72160
rect 32204 72096 32220 72160
rect 32284 72096 32322 72160
rect 31702 72080 32322 72096
rect 31702 72016 31740 72080
rect 31804 72016 31820 72080
rect 31884 72016 31900 72080
rect 31964 72016 31980 72080
rect 32044 72016 32060 72080
rect 32124 72016 32140 72080
rect 32204 72016 32220 72080
rect 32284 72016 32322 72080
rect 31702 72000 32322 72016
rect 31702 71936 31740 72000
rect 31804 71936 31820 72000
rect 31884 71936 31900 72000
rect 31964 71936 31980 72000
rect 32044 71936 32060 72000
rect 32124 71936 32140 72000
rect 32204 71936 32220 72000
rect 32284 71936 32322 72000
rect 31702 62240 32322 71936
rect 31702 62176 31740 62240
rect 31804 62176 31820 62240
rect 31884 62176 31900 62240
rect 31964 62176 31980 62240
rect 32044 62176 32060 62240
rect 32124 62176 32140 62240
rect 32204 62176 32220 62240
rect 32284 62176 32322 62240
rect 31702 62160 32322 62176
rect 31702 62096 31740 62160
rect 31804 62096 31820 62160
rect 31884 62096 31900 62160
rect 31964 62096 31980 62160
rect 32044 62096 32060 62160
rect 32124 62096 32140 62160
rect 32204 62096 32220 62160
rect 32284 62096 32322 62160
rect 31702 62080 32322 62096
rect 31702 62016 31740 62080
rect 31804 62016 31820 62080
rect 31884 62016 31900 62080
rect 31964 62016 31980 62080
rect 32044 62016 32060 62080
rect 32124 62016 32140 62080
rect 32204 62016 32220 62080
rect 32284 62016 32322 62080
rect 31702 62000 32322 62016
rect 31702 61936 31740 62000
rect 31804 61936 31820 62000
rect 31884 61936 31900 62000
rect 31964 61936 31980 62000
rect 32044 61936 32060 62000
rect 32124 61936 32140 62000
rect 32204 61936 32220 62000
rect 32284 61936 32322 62000
rect 31702 52240 32322 61936
rect 31702 52176 31740 52240
rect 31804 52176 31820 52240
rect 31884 52176 31900 52240
rect 31964 52176 31980 52240
rect 32044 52176 32060 52240
rect 32124 52176 32140 52240
rect 32204 52176 32220 52240
rect 32284 52176 32322 52240
rect 31702 52160 32322 52176
rect 31702 52096 31740 52160
rect 31804 52096 31820 52160
rect 31884 52096 31900 52160
rect 31964 52096 31980 52160
rect 32044 52096 32060 52160
rect 32124 52096 32140 52160
rect 32204 52096 32220 52160
rect 32284 52096 32322 52160
rect 31702 52080 32322 52096
rect 31702 52016 31740 52080
rect 31804 52016 31820 52080
rect 31884 52016 31900 52080
rect 31964 52016 31980 52080
rect 32044 52016 32060 52080
rect 32124 52016 32140 52080
rect 32204 52016 32220 52080
rect 32284 52016 32322 52080
rect 31702 52000 32322 52016
rect 31702 51936 31740 52000
rect 31804 51936 31820 52000
rect 31884 51936 31900 52000
rect 31964 51936 31980 52000
rect 32044 51936 32060 52000
rect 32124 51936 32140 52000
rect 32204 51936 32220 52000
rect 32284 51936 32322 52000
rect 31702 42240 32322 51936
rect 31702 42176 31740 42240
rect 31804 42176 31820 42240
rect 31884 42176 31900 42240
rect 31964 42176 31980 42240
rect 32044 42176 32060 42240
rect 32124 42176 32140 42240
rect 32204 42176 32220 42240
rect 32284 42176 32322 42240
rect 31702 42160 32322 42176
rect 31702 42096 31740 42160
rect 31804 42096 31820 42160
rect 31884 42096 31900 42160
rect 31964 42096 31980 42160
rect 32044 42096 32060 42160
rect 32124 42096 32140 42160
rect 32204 42096 32220 42160
rect 32284 42096 32322 42160
rect 31702 42080 32322 42096
rect 31702 42016 31740 42080
rect 31804 42016 31820 42080
rect 31884 42016 31900 42080
rect 31964 42016 31980 42080
rect 32044 42016 32060 42080
rect 32124 42016 32140 42080
rect 32204 42016 32220 42080
rect 32284 42016 32322 42080
rect 31702 42000 32322 42016
rect 31702 41936 31740 42000
rect 31804 41936 31820 42000
rect 31884 41936 31900 42000
rect 31964 41936 31980 42000
rect 32044 41936 32060 42000
rect 32124 41936 32140 42000
rect 32204 41936 32220 42000
rect 32284 41936 32322 42000
rect 31702 32240 32322 41936
rect 31702 32176 31740 32240
rect 31804 32176 31820 32240
rect 31884 32176 31900 32240
rect 31964 32176 31980 32240
rect 32044 32176 32060 32240
rect 32124 32176 32140 32240
rect 32204 32176 32220 32240
rect 32284 32176 32322 32240
rect 31702 32160 32322 32176
rect 31702 32096 31740 32160
rect 31804 32096 31820 32160
rect 31884 32096 31900 32160
rect 31964 32096 31980 32160
rect 32044 32096 32060 32160
rect 32124 32096 32140 32160
rect 32204 32096 32220 32160
rect 32284 32096 32322 32160
rect 31702 32080 32322 32096
rect 31702 32016 31740 32080
rect 31804 32016 31820 32080
rect 31884 32016 31900 32080
rect 31964 32016 31980 32080
rect 32044 32016 32060 32080
rect 32124 32016 32140 32080
rect 32204 32016 32220 32080
rect 32284 32016 32322 32080
rect 31702 32000 32322 32016
rect 31702 31936 31740 32000
rect 31804 31936 31820 32000
rect 31884 31936 31900 32000
rect 31964 31936 31980 32000
rect 32044 31936 32060 32000
rect 32124 31936 32140 32000
rect 32204 31936 32220 32000
rect 32284 31936 32322 32000
rect 31702 22240 32322 31936
rect 31702 22176 31740 22240
rect 31804 22176 31820 22240
rect 31884 22176 31900 22240
rect 31964 22176 31980 22240
rect 32044 22176 32060 22240
rect 32124 22176 32140 22240
rect 32204 22176 32220 22240
rect 32284 22176 32322 22240
rect 31702 22160 32322 22176
rect 31702 22096 31740 22160
rect 31804 22096 31820 22160
rect 31884 22096 31900 22160
rect 31964 22096 31980 22160
rect 32044 22096 32060 22160
rect 32124 22096 32140 22160
rect 32204 22096 32220 22160
rect 32284 22096 32322 22160
rect 31702 22080 32322 22096
rect 31702 22016 31740 22080
rect 31804 22016 31820 22080
rect 31884 22016 31900 22080
rect 31964 22016 31980 22080
rect 32044 22016 32060 22080
rect 32124 22016 32140 22080
rect 32204 22016 32220 22080
rect 32284 22016 32322 22080
rect 31702 22000 32322 22016
rect 31702 21936 31740 22000
rect 31804 21936 31820 22000
rect 31884 21936 31900 22000
rect 31964 21936 31980 22000
rect 32044 21936 32060 22000
rect 32124 21936 32140 22000
rect 32204 21936 32220 22000
rect 32284 21936 32322 22000
rect 31702 12240 32322 21936
rect 31702 12176 31740 12240
rect 31804 12176 31820 12240
rect 31884 12176 31900 12240
rect 31964 12176 31980 12240
rect 32044 12176 32060 12240
rect 32124 12176 32140 12240
rect 32204 12176 32220 12240
rect 32284 12176 32322 12240
rect 31702 12160 32322 12176
rect 31702 12096 31740 12160
rect 31804 12096 31820 12160
rect 31884 12096 31900 12160
rect 31964 12096 31980 12160
rect 32044 12096 32060 12160
rect 32124 12096 32140 12160
rect 32204 12096 32220 12160
rect 32284 12096 32322 12160
rect 31702 12080 32322 12096
rect 31702 12016 31740 12080
rect 31804 12016 31820 12080
rect 31884 12016 31900 12080
rect 31964 12016 31980 12080
rect 32044 12016 32060 12080
rect 32124 12016 32140 12080
rect 32204 12016 32220 12080
rect 32284 12016 32322 12080
rect 31702 12000 32322 12016
rect 31702 11936 31740 12000
rect 31804 11936 31820 12000
rect 31884 11936 31900 12000
rect 31964 11936 31980 12000
rect 32044 11936 32060 12000
rect 32124 11936 32140 12000
rect 32204 11936 32220 12000
rect 32284 11936 32322 12000
rect 31702 2240 32322 11936
rect 34702 84592 35322 87000
rect 34702 84528 34740 84592
rect 34804 84528 34820 84592
rect 34884 84528 34900 84592
rect 34964 84528 34980 84592
rect 35044 84528 35060 84592
rect 35124 84528 35140 84592
rect 35204 84528 35220 84592
rect 35284 84528 35322 84592
rect 34702 84512 35322 84528
rect 34702 84448 34740 84512
rect 34804 84448 34820 84512
rect 34884 84448 34900 84512
rect 34964 84448 34980 84512
rect 35044 84448 35060 84512
rect 35124 84448 35140 84512
rect 35204 84448 35220 84512
rect 35284 84448 35322 84512
rect 34702 84432 35322 84448
rect 34702 84368 34740 84432
rect 34804 84368 34820 84432
rect 34884 84368 34900 84432
rect 34964 84368 34980 84432
rect 35044 84368 35060 84432
rect 35124 84368 35140 84432
rect 35204 84368 35220 84432
rect 35284 84368 35322 84432
rect 34702 84352 35322 84368
rect 34702 84288 34740 84352
rect 34804 84288 34820 84352
rect 34884 84288 34900 84352
rect 34964 84288 34980 84352
rect 35044 84288 35060 84352
rect 35124 84288 35140 84352
rect 35204 84288 35220 84352
rect 35284 84288 35322 84352
rect 34702 74592 35322 84288
rect 34702 74528 34740 74592
rect 34804 74528 34820 74592
rect 34884 74528 34900 74592
rect 34964 74528 34980 74592
rect 35044 74528 35060 74592
rect 35124 74528 35140 74592
rect 35204 74528 35220 74592
rect 35284 74528 35322 74592
rect 34702 74512 35322 74528
rect 34702 74448 34740 74512
rect 34804 74448 34820 74512
rect 34884 74448 34900 74512
rect 34964 74448 34980 74512
rect 35044 74448 35060 74512
rect 35124 74448 35140 74512
rect 35204 74448 35220 74512
rect 35284 74448 35322 74512
rect 34702 74432 35322 74448
rect 34702 74368 34740 74432
rect 34804 74368 34820 74432
rect 34884 74368 34900 74432
rect 34964 74368 34980 74432
rect 35044 74368 35060 74432
rect 35124 74368 35140 74432
rect 35204 74368 35220 74432
rect 35284 74368 35322 74432
rect 34702 74352 35322 74368
rect 34702 74288 34740 74352
rect 34804 74288 34820 74352
rect 34884 74288 34900 74352
rect 34964 74288 34980 74352
rect 35044 74288 35060 74352
rect 35124 74288 35140 74352
rect 35204 74288 35220 74352
rect 35284 74288 35322 74352
rect 34702 64592 35322 74288
rect 34702 64528 34740 64592
rect 34804 64528 34820 64592
rect 34884 64528 34900 64592
rect 34964 64528 34980 64592
rect 35044 64528 35060 64592
rect 35124 64528 35140 64592
rect 35204 64528 35220 64592
rect 35284 64528 35322 64592
rect 34702 64512 35322 64528
rect 34702 64448 34740 64512
rect 34804 64448 34820 64512
rect 34884 64448 34900 64512
rect 34964 64448 34980 64512
rect 35044 64448 35060 64512
rect 35124 64448 35140 64512
rect 35204 64448 35220 64512
rect 35284 64448 35322 64512
rect 34702 64432 35322 64448
rect 34702 64368 34740 64432
rect 34804 64368 34820 64432
rect 34884 64368 34900 64432
rect 34964 64368 34980 64432
rect 35044 64368 35060 64432
rect 35124 64368 35140 64432
rect 35204 64368 35220 64432
rect 35284 64368 35322 64432
rect 34702 64352 35322 64368
rect 34702 64288 34740 64352
rect 34804 64288 34820 64352
rect 34884 64288 34900 64352
rect 34964 64288 34980 64352
rect 35044 64288 35060 64352
rect 35124 64288 35140 64352
rect 35204 64288 35220 64352
rect 35284 64288 35322 64352
rect 34702 54592 35322 64288
rect 34702 54528 34740 54592
rect 34804 54528 34820 54592
rect 34884 54528 34900 54592
rect 34964 54528 34980 54592
rect 35044 54528 35060 54592
rect 35124 54528 35140 54592
rect 35204 54528 35220 54592
rect 35284 54528 35322 54592
rect 34702 54512 35322 54528
rect 34702 54448 34740 54512
rect 34804 54448 34820 54512
rect 34884 54448 34900 54512
rect 34964 54448 34980 54512
rect 35044 54448 35060 54512
rect 35124 54448 35140 54512
rect 35204 54448 35220 54512
rect 35284 54448 35322 54512
rect 34702 54432 35322 54448
rect 34702 54368 34740 54432
rect 34804 54368 34820 54432
rect 34884 54368 34900 54432
rect 34964 54368 34980 54432
rect 35044 54368 35060 54432
rect 35124 54368 35140 54432
rect 35204 54368 35220 54432
rect 35284 54368 35322 54432
rect 34702 54352 35322 54368
rect 34702 54288 34740 54352
rect 34804 54288 34820 54352
rect 34884 54288 34900 54352
rect 34964 54288 34980 54352
rect 35044 54288 35060 54352
rect 35124 54288 35140 54352
rect 35204 54288 35220 54352
rect 35284 54288 35322 54352
rect 34702 44592 35322 54288
rect 34702 44528 34740 44592
rect 34804 44528 34820 44592
rect 34884 44528 34900 44592
rect 34964 44528 34980 44592
rect 35044 44528 35060 44592
rect 35124 44528 35140 44592
rect 35204 44528 35220 44592
rect 35284 44528 35322 44592
rect 34702 44512 35322 44528
rect 34702 44448 34740 44512
rect 34804 44448 34820 44512
rect 34884 44448 34900 44512
rect 34964 44448 34980 44512
rect 35044 44448 35060 44512
rect 35124 44448 35140 44512
rect 35204 44448 35220 44512
rect 35284 44448 35322 44512
rect 34702 44432 35322 44448
rect 34702 44368 34740 44432
rect 34804 44368 34820 44432
rect 34884 44368 34900 44432
rect 34964 44368 34980 44432
rect 35044 44368 35060 44432
rect 35124 44368 35140 44432
rect 35204 44368 35220 44432
rect 35284 44368 35322 44432
rect 34702 44352 35322 44368
rect 34702 44288 34740 44352
rect 34804 44288 34820 44352
rect 34884 44288 34900 44352
rect 34964 44288 34980 44352
rect 35044 44288 35060 44352
rect 35124 44288 35140 44352
rect 35204 44288 35220 44352
rect 35284 44288 35322 44352
rect 34702 34592 35322 44288
rect 34702 34528 34740 34592
rect 34804 34528 34820 34592
rect 34884 34528 34900 34592
rect 34964 34528 34980 34592
rect 35044 34528 35060 34592
rect 35124 34528 35140 34592
rect 35204 34528 35220 34592
rect 35284 34528 35322 34592
rect 34702 34512 35322 34528
rect 34702 34448 34740 34512
rect 34804 34448 34820 34512
rect 34884 34448 34900 34512
rect 34964 34448 34980 34512
rect 35044 34448 35060 34512
rect 35124 34448 35140 34512
rect 35204 34448 35220 34512
rect 35284 34448 35322 34512
rect 34702 34432 35322 34448
rect 34702 34368 34740 34432
rect 34804 34368 34820 34432
rect 34884 34368 34900 34432
rect 34964 34368 34980 34432
rect 35044 34368 35060 34432
rect 35124 34368 35140 34432
rect 35204 34368 35220 34432
rect 35284 34368 35322 34432
rect 34702 34352 35322 34368
rect 34702 34288 34740 34352
rect 34804 34288 34820 34352
rect 34884 34288 34900 34352
rect 34964 34288 34980 34352
rect 35044 34288 35060 34352
rect 35124 34288 35140 34352
rect 35204 34288 35220 34352
rect 35284 34288 35322 34352
rect 34702 24592 35322 34288
rect 34702 24528 34740 24592
rect 34804 24528 34820 24592
rect 34884 24528 34900 24592
rect 34964 24528 34980 24592
rect 35044 24528 35060 24592
rect 35124 24528 35140 24592
rect 35204 24528 35220 24592
rect 35284 24528 35322 24592
rect 34702 24512 35322 24528
rect 34702 24448 34740 24512
rect 34804 24448 34820 24512
rect 34884 24448 34900 24512
rect 34964 24448 34980 24512
rect 35044 24448 35060 24512
rect 35124 24448 35140 24512
rect 35204 24448 35220 24512
rect 35284 24448 35322 24512
rect 34702 24432 35322 24448
rect 34702 24368 34740 24432
rect 34804 24368 34820 24432
rect 34884 24368 34900 24432
rect 34964 24368 34980 24432
rect 35044 24368 35060 24432
rect 35124 24368 35140 24432
rect 35204 24368 35220 24432
rect 35284 24368 35322 24432
rect 34702 24352 35322 24368
rect 34702 24288 34740 24352
rect 34804 24288 34820 24352
rect 34884 24288 34900 24352
rect 34964 24288 34980 24352
rect 35044 24288 35060 24352
rect 35124 24288 35140 24352
rect 35204 24288 35220 24352
rect 35284 24288 35322 24352
rect 34702 14592 35322 24288
rect 34702 14528 34740 14592
rect 34804 14528 34820 14592
rect 34884 14528 34900 14592
rect 34964 14528 34980 14592
rect 35044 14528 35060 14592
rect 35124 14528 35140 14592
rect 35204 14528 35220 14592
rect 35284 14528 35322 14592
rect 34702 14512 35322 14528
rect 34702 14448 34740 14512
rect 34804 14448 34820 14512
rect 34884 14448 34900 14512
rect 34964 14448 34980 14512
rect 35044 14448 35060 14512
rect 35124 14448 35140 14512
rect 35204 14448 35220 14512
rect 35284 14448 35322 14512
rect 34702 14432 35322 14448
rect 34702 14368 34740 14432
rect 34804 14368 34820 14432
rect 34884 14368 34900 14432
rect 34964 14368 34980 14432
rect 35044 14368 35060 14432
rect 35124 14368 35140 14432
rect 35204 14368 35220 14432
rect 35284 14368 35322 14432
rect 34702 14352 35322 14368
rect 34702 14288 34740 14352
rect 34804 14288 34820 14352
rect 34884 14288 34900 14352
rect 34964 14288 34980 14352
rect 35044 14288 35060 14352
rect 35124 14288 35140 14352
rect 35204 14288 35220 14352
rect 35284 14288 35322 14352
rect 33915 4860 33981 4861
rect 33915 4796 33916 4860
rect 33980 4796 33981 4860
rect 33915 4795 33981 4796
rect 33918 2549 33978 4795
rect 34702 4592 35322 14288
rect 34702 4528 34740 4592
rect 34804 4528 34820 4592
rect 34884 4528 34900 4592
rect 34964 4528 34980 4592
rect 35044 4528 35060 4592
rect 35124 4528 35140 4592
rect 35204 4528 35220 4592
rect 35284 4528 35322 4592
rect 34702 4512 35322 4528
rect 34702 4448 34740 4512
rect 34804 4448 34820 4512
rect 34884 4448 34900 4512
rect 34964 4448 34980 4512
rect 35044 4448 35060 4512
rect 35124 4448 35140 4512
rect 35204 4448 35220 4512
rect 35284 4448 35322 4512
rect 34702 4432 35322 4448
rect 34702 4368 34740 4432
rect 34804 4368 34820 4432
rect 34884 4368 34900 4432
rect 34964 4368 34980 4432
rect 35044 4368 35060 4432
rect 35124 4368 35140 4432
rect 35204 4368 35220 4432
rect 35284 4368 35322 4432
rect 34702 4352 35322 4368
rect 34702 4288 34740 4352
rect 34804 4288 34820 4352
rect 34884 4288 34900 4352
rect 34964 4288 34980 4352
rect 35044 4288 35060 4352
rect 35124 4288 35140 4352
rect 35204 4288 35220 4352
rect 35284 4288 35322 4352
rect 33915 2548 33981 2549
rect 33915 2484 33916 2548
rect 33980 2484 33981 2548
rect 33915 2483 33981 2484
rect 31702 2176 31740 2240
rect 31804 2176 31820 2240
rect 31884 2176 31900 2240
rect 31964 2176 31980 2240
rect 32044 2176 32060 2240
rect 32124 2176 32140 2240
rect 32204 2176 32220 2240
rect 32284 2176 32322 2240
rect 31702 2160 32322 2176
rect 31702 2096 31740 2160
rect 31804 2096 31820 2160
rect 31884 2096 31900 2160
rect 31964 2096 31980 2160
rect 32044 2096 32060 2160
rect 32124 2096 32140 2160
rect 32204 2096 32220 2160
rect 32284 2096 32322 2160
rect 31702 2080 32322 2096
rect 31702 2016 31740 2080
rect 31804 2016 31820 2080
rect 31884 2016 31900 2080
rect 31964 2016 31980 2080
rect 32044 2016 32060 2080
rect 32124 2016 32140 2080
rect 32204 2016 32220 2080
rect 32284 2016 32322 2080
rect 31702 2000 32322 2016
rect 31702 1936 31740 2000
rect 31804 1936 31820 2000
rect 31884 1936 31900 2000
rect 31964 1936 31980 2000
rect 32044 1936 32060 2000
rect 32124 1936 32140 2000
rect 32204 1936 32220 2000
rect 32284 1936 32322 2000
rect 31702 0 32322 1936
rect 34702 0 35322 4288
rect 37702 82240 38322 87000
rect 37702 82176 37740 82240
rect 37804 82176 37820 82240
rect 37884 82176 37900 82240
rect 37964 82176 37980 82240
rect 38044 82176 38060 82240
rect 38124 82176 38140 82240
rect 38204 82176 38220 82240
rect 38284 82176 38322 82240
rect 37702 82160 38322 82176
rect 37702 82096 37740 82160
rect 37804 82096 37820 82160
rect 37884 82096 37900 82160
rect 37964 82096 37980 82160
rect 38044 82096 38060 82160
rect 38124 82096 38140 82160
rect 38204 82096 38220 82160
rect 38284 82096 38322 82160
rect 37702 82080 38322 82096
rect 37702 82016 37740 82080
rect 37804 82016 37820 82080
rect 37884 82016 37900 82080
rect 37964 82016 37980 82080
rect 38044 82016 38060 82080
rect 38124 82016 38140 82080
rect 38204 82016 38220 82080
rect 38284 82016 38322 82080
rect 37702 82000 38322 82016
rect 37702 81936 37740 82000
rect 37804 81936 37820 82000
rect 37884 81936 37900 82000
rect 37964 81936 37980 82000
rect 38044 81936 38060 82000
rect 38124 81936 38140 82000
rect 38204 81936 38220 82000
rect 38284 81936 38322 82000
rect 37702 72240 38322 81936
rect 37702 72176 37740 72240
rect 37804 72176 37820 72240
rect 37884 72176 37900 72240
rect 37964 72176 37980 72240
rect 38044 72176 38060 72240
rect 38124 72176 38140 72240
rect 38204 72176 38220 72240
rect 38284 72176 38322 72240
rect 37702 72160 38322 72176
rect 37702 72096 37740 72160
rect 37804 72096 37820 72160
rect 37884 72096 37900 72160
rect 37964 72096 37980 72160
rect 38044 72096 38060 72160
rect 38124 72096 38140 72160
rect 38204 72096 38220 72160
rect 38284 72096 38322 72160
rect 37702 72080 38322 72096
rect 37702 72016 37740 72080
rect 37804 72016 37820 72080
rect 37884 72016 37900 72080
rect 37964 72016 37980 72080
rect 38044 72016 38060 72080
rect 38124 72016 38140 72080
rect 38204 72016 38220 72080
rect 38284 72016 38322 72080
rect 37702 72000 38322 72016
rect 37702 71936 37740 72000
rect 37804 71936 37820 72000
rect 37884 71936 37900 72000
rect 37964 71936 37980 72000
rect 38044 71936 38060 72000
rect 38124 71936 38140 72000
rect 38204 71936 38220 72000
rect 38284 71936 38322 72000
rect 37702 62240 38322 71936
rect 37702 62176 37740 62240
rect 37804 62176 37820 62240
rect 37884 62176 37900 62240
rect 37964 62176 37980 62240
rect 38044 62176 38060 62240
rect 38124 62176 38140 62240
rect 38204 62176 38220 62240
rect 38284 62176 38322 62240
rect 37702 62160 38322 62176
rect 37702 62096 37740 62160
rect 37804 62096 37820 62160
rect 37884 62096 37900 62160
rect 37964 62096 37980 62160
rect 38044 62096 38060 62160
rect 38124 62096 38140 62160
rect 38204 62096 38220 62160
rect 38284 62096 38322 62160
rect 37702 62080 38322 62096
rect 37702 62016 37740 62080
rect 37804 62016 37820 62080
rect 37884 62016 37900 62080
rect 37964 62016 37980 62080
rect 38044 62016 38060 62080
rect 38124 62016 38140 62080
rect 38204 62016 38220 62080
rect 38284 62016 38322 62080
rect 37702 62000 38322 62016
rect 37702 61936 37740 62000
rect 37804 61936 37820 62000
rect 37884 61936 37900 62000
rect 37964 61936 37980 62000
rect 38044 61936 38060 62000
rect 38124 61936 38140 62000
rect 38204 61936 38220 62000
rect 38284 61936 38322 62000
rect 37702 52240 38322 61936
rect 37702 52176 37740 52240
rect 37804 52176 37820 52240
rect 37884 52176 37900 52240
rect 37964 52176 37980 52240
rect 38044 52176 38060 52240
rect 38124 52176 38140 52240
rect 38204 52176 38220 52240
rect 38284 52176 38322 52240
rect 37702 52160 38322 52176
rect 37702 52096 37740 52160
rect 37804 52096 37820 52160
rect 37884 52096 37900 52160
rect 37964 52096 37980 52160
rect 38044 52096 38060 52160
rect 38124 52096 38140 52160
rect 38204 52096 38220 52160
rect 38284 52096 38322 52160
rect 37702 52080 38322 52096
rect 37702 52016 37740 52080
rect 37804 52016 37820 52080
rect 37884 52016 37900 52080
rect 37964 52016 37980 52080
rect 38044 52016 38060 52080
rect 38124 52016 38140 52080
rect 38204 52016 38220 52080
rect 38284 52016 38322 52080
rect 37702 52000 38322 52016
rect 37702 51936 37740 52000
rect 37804 51936 37820 52000
rect 37884 51936 37900 52000
rect 37964 51936 37980 52000
rect 38044 51936 38060 52000
rect 38124 51936 38140 52000
rect 38204 51936 38220 52000
rect 38284 51936 38322 52000
rect 37702 42240 38322 51936
rect 37702 42176 37740 42240
rect 37804 42176 37820 42240
rect 37884 42176 37900 42240
rect 37964 42176 37980 42240
rect 38044 42176 38060 42240
rect 38124 42176 38140 42240
rect 38204 42176 38220 42240
rect 38284 42176 38322 42240
rect 37702 42160 38322 42176
rect 37702 42096 37740 42160
rect 37804 42096 37820 42160
rect 37884 42096 37900 42160
rect 37964 42096 37980 42160
rect 38044 42096 38060 42160
rect 38124 42096 38140 42160
rect 38204 42096 38220 42160
rect 38284 42096 38322 42160
rect 37702 42080 38322 42096
rect 37702 42016 37740 42080
rect 37804 42016 37820 42080
rect 37884 42016 37900 42080
rect 37964 42016 37980 42080
rect 38044 42016 38060 42080
rect 38124 42016 38140 42080
rect 38204 42016 38220 42080
rect 38284 42016 38322 42080
rect 37702 42000 38322 42016
rect 37702 41936 37740 42000
rect 37804 41936 37820 42000
rect 37884 41936 37900 42000
rect 37964 41936 37980 42000
rect 38044 41936 38060 42000
rect 38124 41936 38140 42000
rect 38204 41936 38220 42000
rect 38284 41936 38322 42000
rect 37702 32240 38322 41936
rect 37702 32176 37740 32240
rect 37804 32176 37820 32240
rect 37884 32176 37900 32240
rect 37964 32176 37980 32240
rect 38044 32176 38060 32240
rect 38124 32176 38140 32240
rect 38204 32176 38220 32240
rect 38284 32176 38322 32240
rect 37702 32160 38322 32176
rect 37702 32096 37740 32160
rect 37804 32096 37820 32160
rect 37884 32096 37900 32160
rect 37964 32096 37980 32160
rect 38044 32096 38060 32160
rect 38124 32096 38140 32160
rect 38204 32096 38220 32160
rect 38284 32096 38322 32160
rect 37702 32080 38322 32096
rect 37702 32016 37740 32080
rect 37804 32016 37820 32080
rect 37884 32016 37900 32080
rect 37964 32016 37980 32080
rect 38044 32016 38060 32080
rect 38124 32016 38140 32080
rect 38204 32016 38220 32080
rect 38284 32016 38322 32080
rect 37702 32000 38322 32016
rect 37702 31936 37740 32000
rect 37804 31936 37820 32000
rect 37884 31936 37900 32000
rect 37964 31936 37980 32000
rect 38044 31936 38060 32000
rect 38124 31936 38140 32000
rect 38204 31936 38220 32000
rect 38284 31936 38322 32000
rect 37702 22240 38322 31936
rect 37702 22176 37740 22240
rect 37804 22176 37820 22240
rect 37884 22176 37900 22240
rect 37964 22176 37980 22240
rect 38044 22176 38060 22240
rect 38124 22176 38140 22240
rect 38204 22176 38220 22240
rect 38284 22176 38322 22240
rect 37702 22160 38322 22176
rect 37702 22096 37740 22160
rect 37804 22096 37820 22160
rect 37884 22096 37900 22160
rect 37964 22096 37980 22160
rect 38044 22096 38060 22160
rect 38124 22096 38140 22160
rect 38204 22096 38220 22160
rect 38284 22096 38322 22160
rect 37702 22080 38322 22096
rect 37702 22016 37740 22080
rect 37804 22016 37820 22080
rect 37884 22016 37900 22080
rect 37964 22016 37980 22080
rect 38044 22016 38060 22080
rect 38124 22016 38140 22080
rect 38204 22016 38220 22080
rect 38284 22016 38322 22080
rect 37702 22000 38322 22016
rect 37702 21936 37740 22000
rect 37804 21936 37820 22000
rect 37884 21936 37900 22000
rect 37964 21936 37980 22000
rect 38044 21936 38060 22000
rect 38124 21936 38140 22000
rect 38204 21936 38220 22000
rect 38284 21936 38322 22000
rect 37702 12240 38322 21936
rect 37702 12176 37740 12240
rect 37804 12176 37820 12240
rect 37884 12176 37900 12240
rect 37964 12176 37980 12240
rect 38044 12176 38060 12240
rect 38124 12176 38140 12240
rect 38204 12176 38220 12240
rect 38284 12176 38322 12240
rect 37702 12160 38322 12176
rect 37702 12096 37740 12160
rect 37804 12096 37820 12160
rect 37884 12096 37900 12160
rect 37964 12096 37980 12160
rect 38044 12096 38060 12160
rect 38124 12096 38140 12160
rect 38204 12096 38220 12160
rect 38284 12096 38322 12160
rect 37702 12080 38322 12096
rect 37702 12016 37740 12080
rect 37804 12016 37820 12080
rect 37884 12016 37900 12080
rect 37964 12016 37980 12080
rect 38044 12016 38060 12080
rect 38124 12016 38140 12080
rect 38204 12016 38220 12080
rect 38284 12016 38322 12080
rect 37702 12000 38322 12016
rect 37702 11936 37740 12000
rect 37804 11936 37820 12000
rect 37884 11936 37900 12000
rect 37964 11936 37980 12000
rect 38044 11936 38060 12000
rect 38124 11936 38140 12000
rect 38204 11936 38220 12000
rect 38284 11936 38322 12000
rect 37702 2240 38322 11936
rect 37702 2176 37740 2240
rect 37804 2176 37820 2240
rect 37884 2176 37900 2240
rect 37964 2176 37980 2240
rect 38044 2176 38060 2240
rect 38124 2176 38140 2240
rect 38204 2176 38220 2240
rect 38284 2176 38322 2240
rect 37702 2160 38322 2176
rect 37702 2096 37740 2160
rect 37804 2096 37820 2160
rect 37884 2096 37900 2160
rect 37964 2096 37980 2160
rect 38044 2096 38060 2160
rect 38124 2096 38140 2160
rect 38204 2096 38220 2160
rect 38284 2096 38322 2160
rect 37702 2080 38322 2096
rect 37702 2016 37740 2080
rect 37804 2016 37820 2080
rect 37884 2016 37900 2080
rect 37964 2016 37980 2080
rect 38044 2016 38060 2080
rect 38124 2016 38140 2080
rect 38204 2016 38220 2080
rect 38284 2016 38322 2080
rect 37702 2000 38322 2016
rect 37702 1936 37740 2000
rect 37804 1936 37820 2000
rect 37884 1936 37900 2000
rect 37964 1936 37980 2000
rect 38044 1936 38060 2000
rect 38124 1936 38140 2000
rect 38204 1936 38220 2000
rect 38284 1936 38322 2000
rect 37702 0 38322 1936
rect 40702 84592 41322 87000
rect 40702 84528 40740 84592
rect 40804 84528 40820 84592
rect 40884 84528 40900 84592
rect 40964 84528 40980 84592
rect 41044 84528 41060 84592
rect 41124 84528 41140 84592
rect 41204 84528 41220 84592
rect 41284 84528 41322 84592
rect 40702 84512 41322 84528
rect 40702 84448 40740 84512
rect 40804 84448 40820 84512
rect 40884 84448 40900 84512
rect 40964 84448 40980 84512
rect 41044 84448 41060 84512
rect 41124 84448 41140 84512
rect 41204 84448 41220 84512
rect 41284 84448 41322 84512
rect 40702 84432 41322 84448
rect 40702 84368 40740 84432
rect 40804 84368 40820 84432
rect 40884 84368 40900 84432
rect 40964 84368 40980 84432
rect 41044 84368 41060 84432
rect 41124 84368 41140 84432
rect 41204 84368 41220 84432
rect 41284 84368 41322 84432
rect 40702 84352 41322 84368
rect 40702 84288 40740 84352
rect 40804 84288 40820 84352
rect 40884 84288 40900 84352
rect 40964 84288 40980 84352
rect 41044 84288 41060 84352
rect 41124 84288 41140 84352
rect 41204 84288 41220 84352
rect 41284 84288 41322 84352
rect 40702 74592 41322 84288
rect 40702 74528 40740 74592
rect 40804 74528 40820 74592
rect 40884 74528 40900 74592
rect 40964 74528 40980 74592
rect 41044 74528 41060 74592
rect 41124 74528 41140 74592
rect 41204 74528 41220 74592
rect 41284 74528 41322 74592
rect 40702 74512 41322 74528
rect 40702 74448 40740 74512
rect 40804 74448 40820 74512
rect 40884 74448 40900 74512
rect 40964 74448 40980 74512
rect 41044 74448 41060 74512
rect 41124 74448 41140 74512
rect 41204 74448 41220 74512
rect 41284 74448 41322 74512
rect 40702 74432 41322 74448
rect 40702 74368 40740 74432
rect 40804 74368 40820 74432
rect 40884 74368 40900 74432
rect 40964 74368 40980 74432
rect 41044 74368 41060 74432
rect 41124 74368 41140 74432
rect 41204 74368 41220 74432
rect 41284 74368 41322 74432
rect 40702 74352 41322 74368
rect 40702 74288 40740 74352
rect 40804 74288 40820 74352
rect 40884 74288 40900 74352
rect 40964 74288 40980 74352
rect 41044 74288 41060 74352
rect 41124 74288 41140 74352
rect 41204 74288 41220 74352
rect 41284 74288 41322 74352
rect 40702 64592 41322 74288
rect 40702 64528 40740 64592
rect 40804 64528 40820 64592
rect 40884 64528 40900 64592
rect 40964 64528 40980 64592
rect 41044 64528 41060 64592
rect 41124 64528 41140 64592
rect 41204 64528 41220 64592
rect 41284 64528 41322 64592
rect 40702 64512 41322 64528
rect 40702 64448 40740 64512
rect 40804 64448 40820 64512
rect 40884 64448 40900 64512
rect 40964 64448 40980 64512
rect 41044 64448 41060 64512
rect 41124 64448 41140 64512
rect 41204 64448 41220 64512
rect 41284 64448 41322 64512
rect 40702 64432 41322 64448
rect 40702 64368 40740 64432
rect 40804 64368 40820 64432
rect 40884 64368 40900 64432
rect 40964 64368 40980 64432
rect 41044 64368 41060 64432
rect 41124 64368 41140 64432
rect 41204 64368 41220 64432
rect 41284 64368 41322 64432
rect 40702 64352 41322 64368
rect 40702 64288 40740 64352
rect 40804 64288 40820 64352
rect 40884 64288 40900 64352
rect 40964 64288 40980 64352
rect 41044 64288 41060 64352
rect 41124 64288 41140 64352
rect 41204 64288 41220 64352
rect 41284 64288 41322 64352
rect 40702 54592 41322 64288
rect 40702 54528 40740 54592
rect 40804 54528 40820 54592
rect 40884 54528 40900 54592
rect 40964 54528 40980 54592
rect 41044 54528 41060 54592
rect 41124 54528 41140 54592
rect 41204 54528 41220 54592
rect 41284 54528 41322 54592
rect 40702 54512 41322 54528
rect 40702 54448 40740 54512
rect 40804 54448 40820 54512
rect 40884 54448 40900 54512
rect 40964 54448 40980 54512
rect 41044 54448 41060 54512
rect 41124 54448 41140 54512
rect 41204 54448 41220 54512
rect 41284 54448 41322 54512
rect 40702 54432 41322 54448
rect 40702 54368 40740 54432
rect 40804 54368 40820 54432
rect 40884 54368 40900 54432
rect 40964 54368 40980 54432
rect 41044 54368 41060 54432
rect 41124 54368 41140 54432
rect 41204 54368 41220 54432
rect 41284 54368 41322 54432
rect 40702 54352 41322 54368
rect 40702 54288 40740 54352
rect 40804 54288 40820 54352
rect 40884 54288 40900 54352
rect 40964 54288 40980 54352
rect 41044 54288 41060 54352
rect 41124 54288 41140 54352
rect 41204 54288 41220 54352
rect 41284 54288 41322 54352
rect 40702 44592 41322 54288
rect 40702 44528 40740 44592
rect 40804 44528 40820 44592
rect 40884 44528 40900 44592
rect 40964 44528 40980 44592
rect 41044 44528 41060 44592
rect 41124 44528 41140 44592
rect 41204 44528 41220 44592
rect 41284 44528 41322 44592
rect 40702 44512 41322 44528
rect 40702 44448 40740 44512
rect 40804 44448 40820 44512
rect 40884 44448 40900 44512
rect 40964 44448 40980 44512
rect 41044 44448 41060 44512
rect 41124 44448 41140 44512
rect 41204 44448 41220 44512
rect 41284 44448 41322 44512
rect 40702 44432 41322 44448
rect 40702 44368 40740 44432
rect 40804 44368 40820 44432
rect 40884 44368 40900 44432
rect 40964 44368 40980 44432
rect 41044 44368 41060 44432
rect 41124 44368 41140 44432
rect 41204 44368 41220 44432
rect 41284 44368 41322 44432
rect 40702 44352 41322 44368
rect 40702 44288 40740 44352
rect 40804 44288 40820 44352
rect 40884 44288 40900 44352
rect 40964 44288 40980 44352
rect 41044 44288 41060 44352
rect 41124 44288 41140 44352
rect 41204 44288 41220 44352
rect 41284 44288 41322 44352
rect 40702 34592 41322 44288
rect 40702 34528 40740 34592
rect 40804 34528 40820 34592
rect 40884 34528 40900 34592
rect 40964 34528 40980 34592
rect 41044 34528 41060 34592
rect 41124 34528 41140 34592
rect 41204 34528 41220 34592
rect 41284 34528 41322 34592
rect 40702 34512 41322 34528
rect 40702 34448 40740 34512
rect 40804 34448 40820 34512
rect 40884 34448 40900 34512
rect 40964 34448 40980 34512
rect 41044 34448 41060 34512
rect 41124 34448 41140 34512
rect 41204 34448 41220 34512
rect 41284 34448 41322 34512
rect 40702 34432 41322 34448
rect 40702 34368 40740 34432
rect 40804 34368 40820 34432
rect 40884 34368 40900 34432
rect 40964 34368 40980 34432
rect 41044 34368 41060 34432
rect 41124 34368 41140 34432
rect 41204 34368 41220 34432
rect 41284 34368 41322 34432
rect 40702 34352 41322 34368
rect 40702 34288 40740 34352
rect 40804 34288 40820 34352
rect 40884 34288 40900 34352
rect 40964 34288 40980 34352
rect 41044 34288 41060 34352
rect 41124 34288 41140 34352
rect 41204 34288 41220 34352
rect 41284 34288 41322 34352
rect 40702 24592 41322 34288
rect 40702 24528 40740 24592
rect 40804 24528 40820 24592
rect 40884 24528 40900 24592
rect 40964 24528 40980 24592
rect 41044 24528 41060 24592
rect 41124 24528 41140 24592
rect 41204 24528 41220 24592
rect 41284 24528 41322 24592
rect 40702 24512 41322 24528
rect 40702 24448 40740 24512
rect 40804 24448 40820 24512
rect 40884 24448 40900 24512
rect 40964 24448 40980 24512
rect 41044 24448 41060 24512
rect 41124 24448 41140 24512
rect 41204 24448 41220 24512
rect 41284 24448 41322 24512
rect 40702 24432 41322 24448
rect 40702 24368 40740 24432
rect 40804 24368 40820 24432
rect 40884 24368 40900 24432
rect 40964 24368 40980 24432
rect 41044 24368 41060 24432
rect 41124 24368 41140 24432
rect 41204 24368 41220 24432
rect 41284 24368 41322 24432
rect 40702 24352 41322 24368
rect 40702 24288 40740 24352
rect 40804 24288 40820 24352
rect 40884 24288 40900 24352
rect 40964 24288 40980 24352
rect 41044 24288 41060 24352
rect 41124 24288 41140 24352
rect 41204 24288 41220 24352
rect 41284 24288 41322 24352
rect 40702 14592 41322 24288
rect 40702 14528 40740 14592
rect 40804 14528 40820 14592
rect 40884 14528 40900 14592
rect 40964 14528 40980 14592
rect 41044 14528 41060 14592
rect 41124 14528 41140 14592
rect 41204 14528 41220 14592
rect 41284 14528 41322 14592
rect 40702 14512 41322 14528
rect 40702 14448 40740 14512
rect 40804 14448 40820 14512
rect 40884 14448 40900 14512
rect 40964 14448 40980 14512
rect 41044 14448 41060 14512
rect 41124 14448 41140 14512
rect 41204 14448 41220 14512
rect 41284 14448 41322 14512
rect 40702 14432 41322 14448
rect 40702 14368 40740 14432
rect 40804 14368 40820 14432
rect 40884 14368 40900 14432
rect 40964 14368 40980 14432
rect 41044 14368 41060 14432
rect 41124 14368 41140 14432
rect 41204 14368 41220 14432
rect 41284 14368 41322 14432
rect 40702 14352 41322 14368
rect 40702 14288 40740 14352
rect 40804 14288 40820 14352
rect 40884 14288 40900 14352
rect 40964 14288 40980 14352
rect 41044 14288 41060 14352
rect 41124 14288 41140 14352
rect 41204 14288 41220 14352
rect 41284 14288 41322 14352
rect 40702 4592 41322 14288
rect 40702 4528 40740 4592
rect 40804 4528 40820 4592
rect 40884 4528 40900 4592
rect 40964 4528 40980 4592
rect 41044 4528 41060 4592
rect 41124 4528 41140 4592
rect 41204 4528 41220 4592
rect 41284 4528 41322 4592
rect 40702 4512 41322 4528
rect 40702 4448 40740 4512
rect 40804 4448 40820 4512
rect 40884 4448 40900 4512
rect 40964 4448 40980 4512
rect 41044 4448 41060 4512
rect 41124 4448 41140 4512
rect 41204 4448 41220 4512
rect 41284 4448 41322 4512
rect 40702 4432 41322 4448
rect 40702 4368 40740 4432
rect 40804 4368 40820 4432
rect 40884 4368 40900 4432
rect 40964 4368 40980 4432
rect 41044 4368 41060 4432
rect 41124 4368 41140 4432
rect 41204 4368 41220 4432
rect 41284 4368 41322 4432
rect 40702 4352 41322 4368
rect 40702 4288 40740 4352
rect 40804 4288 40820 4352
rect 40884 4288 40900 4352
rect 40964 4288 40980 4352
rect 41044 4288 41060 4352
rect 41124 4288 41140 4352
rect 41204 4288 41220 4352
rect 41284 4288 41322 4352
rect 40702 0 41322 4288
rect 43702 82240 44322 87000
rect 43702 82176 43740 82240
rect 43804 82176 43820 82240
rect 43884 82176 43900 82240
rect 43964 82176 43980 82240
rect 44044 82176 44060 82240
rect 44124 82176 44140 82240
rect 44204 82176 44220 82240
rect 44284 82176 44322 82240
rect 43702 82160 44322 82176
rect 43702 82096 43740 82160
rect 43804 82096 43820 82160
rect 43884 82096 43900 82160
rect 43964 82096 43980 82160
rect 44044 82096 44060 82160
rect 44124 82096 44140 82160
rect 44204 82096 44220 82160
rect 44284 82096 44322 82160
rect 43702 82080 44322 82096
rect 43702 82016 43740 82080
rect 43804 82016 43820 82080
rect 43884 82016 43900 82080
rect 43964 82016 43980 82080
rect 44044 82016 44060 82080
rect 44124 82016 44140 82080
rect 44204 82016 44220 82080
rect 44284 82016 44322 82080
rect 43702 82000 44322 82016
rect 43702 81936 43740 82000
rect 43804 81936 43820 82000
rect 43884 81936 43900 82000
rect 43964 81936 43980 82000
rect 44044 81936 44060 82000
rect 44124 81936 44140 82000
rect 44204 81936 44220 82000
rect 44284 81936 44322 82000
rect 43702 72240 44322 81936
rect 43702 72176 43740 72240
rect 43804 72176 43820 72240
rect 43884 72176 43900 72240
rect 43964 72176 43980 72240
rect 44044 72176 44060 72240
rect 44124 72176 44140 72240
rect 44204 72176 44220 72240
rect 44284 72176 44322 72240
rect 43702 72160 44322 72176
rect 43702 72096 43740 72160
rect 43804 72096 43820 72160
rect 43884 72096 43900 72160
rect 43964 72096 43980 72160
rect 44044 72096 44060 72160
rect 44124 72096 44140 72160
rect 44204 72096 44220 72160
rect 44284 72096 44322 72160
rect 43702 72080 44322 72096
rect 43702 72016 43740 72080
rect 43804 72016 43820 72080
rect 43884 72016 43900 72080
rect 43964 72016 43980 72080
rect 44044 72016 44060 72080
rect 44124 72016 44140 72080
rect 44204 72016 44220 72080
rect 44284 72016 44322 72080
rect 43702 72000 44322 72016
rect 43702 71936 43740 72000
rect 43804 71936 43820 72000
rect 43884 71936 43900 72000
rect 43964 71936 43980 72000
rect 44044 71936 44060 72000
rect 44124 71936 44140 72000
rect 44204 71936 44220 72000
rect 44284 71936 44322 72000
rect 43702 62240 44322 71936
rect 43702 62176 43740 62240
rect 43804 62176 43820 62240
rect 43884 62176 43900 62240
rect 43964 62176 43980 62240
rect 44044 62176 44060 62240
rect 44124 62176 44140 62240
rect 44204 62176 44220 62240
rect 44284 62176 44322 62240
rect 43702 62160 44322 62176
rect 43702 62096 43740 62160
rect 43804 62096 43820 62160
rect 43884 62096 43900 62160
rect 43964 62096 43980 62160
rect 44044 62096 44060 62160
rect 44124 62096 44140 62160
rect 44204 62096 44220 62160
rect 44284 62096 44322 62160
rect 43702 62080 44322 62096
rect 43702 62016 43740 62080
rect 43804 62016 43820 62080
rect 43884 62016 43900 62080
rect 43964 62016 43980 62080
rect 44044 62016 44060 62080
rect 44124 62016 44140 62080
rect 44204 62016 44220 62080
rect 44284 62016 44322 62080
rect 43702 62000 44322 62016
rect 43702 61936 43740 62000
rect 43804 61936 43820 62000
rect 43884 61936 43900 62000
rect 43964 61936 43980 62000
rect 44044 61936 44060 62000
rect 44124 61936 44140 62000
rect 44204 61936 44220 62000
rect 44284 61936 44322 62000
rect 43702 52240 44322 61936
rect 43702 52176 43740 52240
rect 43804 52176 43820 52240
rect 43884 52176 43900 52240
rect 43964 52176 43980 52240
rect 44044 52176 44060 52240
rect 44124 52176 44140 52240
rect 44204 52176 44220 52240
rect 44284 52176 44322 52240
rect 43702 52160 44322 52176
rect 43702 52096 43740 52160
rect 43804 52096 43820 52160
rect 43884 52096 43900 52160
rect 43964 52096 43980 52160
rect 44044 52096 44060 52160
rect 44124 52096 44140 52160
rect 44204 52096 44220 52160
rect 44284 52096 44322 52160
rect 43702 52080 44322 52096
rect 43702 52016 43740 52080
rect 43804 52016 43820 52080
rect 43884 52016 43900 52080
rect 43964 52016 43980 52080
rect 44044 52016 44060 52080
rect 44124 52016 44140 52080
rect 44204 52016 44220 52080
rect 44284 52016 44322 52080
rect 43702 52000 44322 52016
rect 43702 51936 43740 52000
rect 43804 51936 43820 52000
rect 43884 51936 43900 52000
rect 43964 51936 43980 52000
rect 44044 51936 44060 52000
rect 44124 51936 44140 52000
rect 44204 51936 44220 52000
rect 44284 51936 44322 52000
rect 43702 42240 44322 51936
rect 43702 42176 43740 42240
rect 43804 42176 43820 42240
rect 43884 42176 43900 42240
rect 43964 42176 43980 42240
rect 44044 42176 44060 42240
rect 44124 42176 44140 42240
rect 44204 42176 44220 42240
rect 44284 42176 44322 42240
rect 43702 42160 44322 42176
rect 43702 42096 43740 42160
rect 43804 42096 43820 42160
rect 43884 42096 43900 42160
rect 43964 42096 43980 42160
rect 44044 42096 44060 42160
rect 44124 42096 44140 42160
rect 44204 42096 44220 42160
rect 44284 42096 44322 42160
rect 43702 42080 44322 42096
rect 43702 42016 43740 42080
rect 43804 42016 43820 42080
rect 43884 42016 43900 42080
rect 43964 42016 43980 42080
rect 44044 42016 44060 42080
rect 44124 42016 44140 42080
rect 44204 42016 44220 42080
rect 44284 42016 44322 42080
rect 43702 42000 44322 42016
rect 43702 41936 43740 42000
rect 43804 41936 43820 42000
rect 43884 41936 43900 42000
rect 43964 41936 43980 42000
rect 44044 41936 44060 42000
rect 44124 41936 44140 42000
rect 44204 41936 44220 42000
rect 44284 41936 44322 42000
rect 43702 32240 44322 41936
rect 43702 32176 43740 32240
rect 43804 32176 43820 32240
rect 43884 32176 43900 32240
rect 43964 32176 43980 32240
rect 44044 32176 44060 32240
rect 44124 32176 44140 32240
rect 44204 32176 44220 32240
rect 44284 32176 44322 32240
rect 43702 32160 44322 32176
rect 43702 32096 43740 32160
rect 43804 32096 43820 32160
rect 43884 32096 43900 32160
rect 43964 32096 43980 32160
rect 44044 32096 44060 32160
rect 44124 32096 44140 32160
rect 44204 32096 44220 32160
rect 44284 32096 44322 32160
rect 43702 32080 44322 32096
rect 43702 32016 43740 32080
rect 43804 32016 43820 32080
rect 43884 32016 43900 32080
rect 43964 32016 43980 32080
rect 44044 32016 44060 32080
rect 44124 32016 44140 32080
rect 44204 32016 44220 32080
rect 44284 32016 44322 32080
rect 43702 32000 44322 32016
rect 43702 31936 43740 32000
rect 43804 31936 43820 32000
rect 43884 31936 43900 32000
rect 43964 31936 43980 32000
rect 44044 31936 44060 32000
rect 44124 31936 44140 32000
rect 44204 31936 44220 32000
rect 44284 31936 44322 32000
rect 43702 22240 44322 31936
rect 43702 22176 43740 22240
rect 43804 22176 43820 22240
rect 43884 22176 43900 22240
rect 43964 22176 43980 22240
rect 44044 22176 44060 22240
rect 44124 22176 44140 22240
rect 44204 22176 44220 22240
rect 44284 22176 44322 22240
rect 43702 22160 44322 22176
rect 43702 22096 43740 22160
rect 43804 22096 43820 22160
rect 43884 22096 43900 22160
rect 43964 22096 43980 22160
rect 44044 22096 44060 22160
rect 44124 22096 44140 22160
rect 44204 22096 44220 22160
rect 44284 22096 44322 22160
rect 43702 22080 44322 22096
rect 43702 22016 43740 22080
rect 43804 22016 43820 22080
rect 43884 22016 43900 22080
rect 43964 22016 43980 22080
rect 44044 22016 44060 22080
rect 44124 22016 44140 22080
rect 44204 22016 44220 22080
rect 44284 22016 44322 22080
rect 43702 22000 44322 22016
rect 43702 21936 43740 22000
rect 43804 21936 43820 22000
rect 43884 21936 43900 22000
rect 43964 21936 43980 22000
rect 44044 21936 44060 22000
rect 44124 21936 44140 22000
rect 44204 21936 44220 22000
rect 44284 21936 44322 22000
rect 43702 12240 44322 21936
rect 43702 12176 43740 12240
rect 43804 12176 43820 12240
rect 43884 12176 43900 12240
rect 43964 12176 43980 12240
rect 44044 12176 44060 12240
rect 44124 12176 44140 12240
rect 44204 12176 44220 12240
rect 44284 12176 44322 12240
rect 43702 12160 44322 12176
rect 43702 12096 43740 12160
rect 43804 12096 43820 12160
rect 43884 12096 43900 12160
rect 43964 12096 43980 12160
rect 44044 12096 44060 12160
rect 44124 12096 44140 12160
rect 44204 12096 44220 12160
rect 44284 12096 44322 12160
rect 43702 12080 44322 12096
rect 43702 12016 43740 12080
rect 43804 12016 43820 12080
rect 43884 12016 43900 12080
rect 43964 12016 43980 12080
rect 44044 12016 44060 12080
rect 44124 12016 44140 12080
rect 44204 12016 44220 12080
rect 44284 12016 44322 12080
rect 43702 12000 44322 12016
rect 43702 11936 43740 12000
rect 43804 11936 43820 12000
rect 43884 11936 43900 12000
rect 43964 11936 43980 12000
rect 44044 11936 44060 12000
rect 44124 11936 44140 12000
rect 44204 11936 44220 12000
rect 44284 11936 44322 12000
rect 43702 2240 44322 11936
rect 43702 2176 43740 2240
rect 43804 2176 43820 2240
rect 43884 2176 43900 2240
rect 43964 2176 43980 2240
rect 44044 2176 44060 2240
rect 44124 2176 44140 2240
rect 44204 2176 44220 2240
rect 44284 2176 44322 2240
rect 43702 2160 44322 2176
rect 43702 2096 43740 2160
rect 43804 2096 43820 2160
rect 43884 2096 43900 2160
rect 43964 2096 43980 2160
rect 44044 2096 44060 2160
rect 44124 2096 44140 2160
rect 44204 2096 44220 2160
rect 44284 2096 44322 2160
rect 43702 2080 44322 2096
rect 43702 2016 43740 2080
rect 43804 2016 43820 2080
rect 43884 2016 43900 2080
rect 43964 2016 43980 2080
rect 44044 2016 44060 2080
rect 44124 2016 44140 2080
rect 44204 2016 44220 2080
rect 44284 2016 44322 2080
rect 43702 2000 44322 2016
rect 43702 1936 43740 2000
rect 43804 1936 43820 2000
rect 43884 1936 43900 2000
rect 43964 1936 43980 2000
rect 44044 1936 44060 2000
rect 44124 1936 44140 2000
rect 44204 1936 44220 2000
rect 44284 1936 44322 2000
rect 43702 0 44322 1936
rect 46702 84592 47322 87000
rect 46702 84528 46740 84592
rect 46804 84528 46820 84592
rect 46884 84528 46900 84592
rect 46964 84528 46980 84592
rect 47044 84528 47060 84592
rect 47124 84528 47140 84592
rect 47204 84528 47220 84592
rect 47284 84528 47322 84592
rect 46702 84512 47322 84528
rect 46702 84448 46740 84512
rect 46804 84448 46820 84512
rect 46884 84448 46900 84512
rect 46964 84448 46980 84512
rect 47044 84448 47060 84512
rect 47124 84448 47140 84512
rect 47204 84448 47220 84512
rect 47284 84448 47322 84512
rect 46702 84432 47322 84448
rect 46702 84368 46740 84432
rect 46804 84368 46820 84432
rect 46884 84368 46900 84432
rect 46964 84368 46980 84432
rect 47044 84368 47060 84432
rect 47124 84368 47140 84432
rect 47204 84368 47220 84432
rect 47284 84368 47322 84432
rect 46702 84352 47322 84368
rect 46702 84288 46740 84352
rect 46804 84288 46820 84352
rect 46884 84288 46900 84352
rect 46964 84288 46980 84352
rect 47044 84288 47060 84352
rect 47124 84288 47140 84352
rect 47204 84288 47220 84352
rect 47284 84288 47322 84352
rect 46702 74592 47322 84288
rect 46702 74528 46740 74592
rect 46804 74528 46820 74592
rect 46884 74528 46900 74592
rect 46964 74528 46980 74592
rect 47044 74528 47060 74592
rect 47124 74528 47140 74592
rect 47204 74528 47220 74592
rect 47284 74528 47322 74592
rect 46702 74512 47322 74528
rect 46702 74448 46740 74512
rect 46804 74448 46820 74512
rect 46884 74448 46900 74512
rect 46964 74448 46980 74512
rect 47044 74448 47060 74512
rect 47124 74448 47140 74512
rect 47204 74448 47220 74512
rect 47284 74448 47322 74512
rect 46702 74432 47322 74448
rect 46702 74368 46740 74432
rect 46804 74368 46820 74432
rect 46884 74368 46900 74432
rect 46964 74368 46980 74432
rect 47044 74368 47060 74432
rect 47124 74368 47140 74432
rect 47204 74368 47220 74432
rect 47284 74368 47322 74432
rect 46702 74352 47322 74368
rect 46702 74288 46740 74352
rect 46804 74288 46820 74352
rect 46884 74288 46900 74352
rect 46964 74288 46980 74352
rect 47044 74288 47060 74352
rect 47124 74288 47140 74352
rect 47204 74288 47220 74352
rect 47284 74288 47322 74352
rect 46702 64592 47322 74288
rect 46702 64528 46740 64592
rect 46804 64528 46820 64592
rect 46884 64528 46900 64592
rect 46964 64528 46980 64592
rect 47044 64528 47060 64592
rect 47124 64528 47140 64592
rect 47204 64528 47220 64592
rect 47284 64528 47322 64592
rect 46702 64512 47322 64528
rect 46702 64448 46740 64512
rect 46804 64448 46820 64512
rect 46884 64448 46900 64512
rect 46964 64448 46980 64512
rect 47044 64448 47060 64512
rect 47124 64448 47140 64512
rect 47204 64448 47220 64512
rect 47284 64448 47322 64512
rect 46702 64432 47322 64448
rect 46702 64368 46740 64432
rect 46804 64368 46820 64432
rect 46884 64368 46900 64432
rect 46964 64368 46980 64432
rect 47044 64368 47060 64432
rect 47124 64368 47140 64432
rect 47204 64368 47220 64432
rect 47284 64368 47322 64432
rect 46702 64352 47322 64368
rect 46702 64288 46740 64352
rect 46804 64288 46820 64352
rect 46884 64288 46900 64352
rect 46964 64288 46980 64352
rect 47044 64288 47060 64352
rect 47124 64288 47140 64352
rect 47204 64288 47220 64352
rect 47284 64288 47322 64352
rect 46702 54592 47322 64288
rect 46702 54528 46740 54592
rect 46804 54528 46820 54592
rect 46884 54528 46900 54592
rect 46964 54528 46980 54592
rect 47044 54528 47060 54592
rect 47124 54528 47140 54592
rect 47204 54528 47220 54592
rect 47284 54528 47322 54592
rect 46702 54512 47322 54528
rect 46702 54448 46740 54512
rect 46804 54448 46820 54512
rect 46884 54448 46900 54512
rect 46964 54448 46980 54512
rect 47044 54448 47060 54512
rect 47124 54448 47140 54512
rect 47204 54448 47220 54512
rect 47284 54448 47322 54512
rect 46702 54432 47322 54448
rect 46702 54368 46740 54432
rect 46804 54368 46820 54432
rect 46884 54368 46900 54432
rect 46964 54368 46980 54432
rect 47044 54368 47060 54432
rect 47124 54368 47140 54432
rect 47204 54368 47220 54432
rect 47284 54368 47322 54432
rect 46702 54352 47322 54368
rect 46702 54288 46740 54352
rect 46804 54288 46820 54352
rect 46884 54288 46900 54352
rect 46964 54288 46980 54352
rect 47044 54288 47060 54352
rect 47124 54288 47140 54352
rect 47204 54288 47220 54352
rect 47284 54288 47322 54352
rect 46702 44592 47322 54288
rect 46702 44528 46740 44592
rect 46804 44528 46820 44592
rect 46884 44528 46900 44592
rect 46964 44528 46980 44592
rect 47044 44528 47060 44592
rect 47124 44528 47140 44592
rect 47204 44528 47220 44592
rect 47284 44528 47322 44592
rect 46702 44512 47322 44528
rect 46702 44448 46740 44512
rect 46804 44448 46820 44512
rect 46884 44448 46900 44512
rect 46964 44448 46980 44512
rect 47044 44448 47060 44512
rect 47124 44448 47140 44512
rect 47204 44448 47220 44512
rect 47284 44448 47322 44512
rect 46702 44432 47322 44448
rect 46702 44368 46740 44432
rect 46804 44368 46820 44432
rect 46884 44368 46900 44432
rect 46964 44368 46980 44432
rect 47044 44368 47060 44432
rect 47124 44368 47140 44432
rect 47204 44368 47220 44432
rect 47284 44368 47322 44432
rect 46702 44352 47322 44368
rect 46702 44288 46740 44352
rect 46804 44288 46820 44352
rect 46884 44288 46900 44352
rect 46964 44288 46980 44352
rect 47044 44288 47060 44352
rect 47124 44288 47140 44352
rect 47204 44288 47220 44352
rect 47284 44288 47322 44352
rect 46702 34592 47322 44288
rect 46702 34528 46740 34592
rect 46804 34528 46820 34592
rect 46884 34528 46900 34592
rect 46964 34528 46980 34592
rect 47044 34528 47060 34592
rect 47124 34528 47140 34592
rect 47204 34528 47220 34592
rect 47284 34528 47322 34592
rect 46702 34512 47322 34528
rect 46702 34448 46740 34512
rect 46804 34448 46820 34512
rect 46884 34448 46900 34512
rect 46964 34448 46980 34512
rect 47044 34448 47060 34512
rect 47124 34448 47140 34512
rect 47204 34448 47220 34512
rect 47284 34448 47322 34512
rect 46702 34432 47322 34448
rect 46702 34368 46740 34432
rect 46804 34368 46820 34432
rect 46884 34368 46900 34432
rect 46964 34368 46980 34432
rect 47044 34368 47060 34432
rect 47124 34368 47140 34432
rect 47204 34368 47220 34432
rect 47284 34368 47322 34432
rect 46702 34352 47322 34368
rect 46702 34288 46740 34352
rect 46804 34288 46820 34352
rect 46884 34288 46900 34352
rect 46964 34288 46980 34352
rect 47044 34288 47060 34352
rect 47124 34288 47140 34352
rect 47204 34288 47220 34352
rect 47284 34288 47322 34352
rect 46702 24592 47322 34288
rect 46702 24528 46740 24592
rect 46804 24528 46820 24592
rect 46884 24528 46900 24592
rect 46964 24528 46980 24592
rect 47044 24528 47060 24592
rect 47124 24528 47140 24592
rect 47204 24528 47220 24592
rect 47284 24528 47322 24592
rect 46702 24512 47322 24528
rect 46702 24448 46740 24512
rect 46804 24448 46820 24512
rect 46884 24448 46900 24512
rect 46964 24448 46980 24512
rect 47044 24448 47060 24512
rect 47124 24448 47140 24512
rect 47204 24448 47220 24512
rect 47284 24448 47322 24512
rect 46702 24432 47322 24448
rect 46702 24368 46740 24432
rect 46804 24368 46820 24432
rect 46884 24368 46900 24432
rect 46964 24368 46980 24432
rect 47044 24368 47060 24432
rect 47124 24368 47140 24432
rect 47204 24368 47220 24432
rect 47284 24368 47322 24432
rect 46702 24352 47322 24368
rect 46702 24288 46740 24352
rect 46804 24288 46820 24352
rect 46884 24288 46900 24352
rect 46964 24288 46980 24352
rect 47044 24288 47060 24352
rect 47124 24288 47140 24352
rect 47204 24288 47220 24352
rect 47284 24288 47322 24352
rect 46702 14592 47322 24288
rect 46702 14528 46740 14592
rect 46804 14528 46820 14592
rect 46884 14528 46900 14592
rect 46964 14528 46980 14592
rect 47044 14528 47060 14592
rect 47124 14528 47140 14592
rect 47204 14528 47220 14592
rect 47284 14528 47322 14592
rect 46702 14512 47322 14528
rect 46702 14448 46740 14512
rect 46804 14448 46820 14512
rect 46884 14448 46900 14512
rect 46964 14448 46980 14512
rect 47044 14448 47060 14512
rect 47124 14448 47140 14512
rect 47204 14448 47220 14512
rect 47284 14448 47322 14512
rect 46702 14432 47322 14448
rect 46702 14368 46740 14432
rect 46804 14368 46820 14432
rect 46884 14368 46900 14432
rect 46964 14368 46980 14432
rect 47044 14368 47060 14432
rect 47124 14368 47140 14432
rect 47204 14368 47220 14432
rect 47284 14368 47322 14432
rect 46702 14352 47322 14368
rect 46702 14288 46740 14352
rect 46804 14288 46820 14352
rect 46884 14288 46900 14352
rect 46964 14288 46980 14352
rect 47044 14288 47060 14352
rect 47124 14288 47140 14352
rect 47204 14288 47220 14352
rect 47284 14288 47322 14352
rect 46702 4592 47322 14288
rect 46702 4528 46740 4592
rect 46804 4528 46820 4592
rect 46884 4528 46900 4592
rect 46964 4528 46980 4592
rect 47044 4528 47060 4592
rect 47124 4528 47140 4592
rect 47204 4528 47220 4592
rect 47284 4528 47322 4592
rect 46702 4512 47322 4528
rect 46702 4448 46740 4512
rect 46804 4448 46820 4512
rect 46884 4448 46900 4512
rect 46964 4448 46980 4512
rect 47044 4448 47060 4512
rect 47124 4448 47140 4512
rect 47204 4448 47220 4512
rect 47284 4448 47322 4512
rect 46702 4432 47322 4448
rect 46702 4368 46740 4432
rect 46804 4368 46820 4432
rect 46884 4368 46900 4432
rect 46964 4368 46980 4432
rect 47044 4368 47060 4432
rect 47124 4368 47140 4432
rect 47204 4368 47220 4432
rect 47284 4368 47322 4432
rect 46702 4352 47322 4368
rect 46702 4288 46740 4352
rect 46804 4288 46820 4352
rect 46884 4288 46900 4352
rect 46964 4288 46980 4352
rect 47044 4288 47060 4352
rect 47124 4288 47140 4352
rect 47204 4288 47220 4352
rect 47284 4288 47322 4352
rect 46702 0 47322 4288
rect 49702 82240 50322 87000
rect 49702 82176 49740 82240
rect 49804 82176 49820 82240
rect 49884 82176 49900 82240
rect 49964 82176 49980 82240
rect 50044 82176 50060 82240
rect 50124 82176 50140 82240
rect 50204 82176 50220 82240
rect 50284 82176 50322 82240
rect 49702 82160 50322 82176
rect 49702 82096 49740 82160
rect 49804 82096 49820 82160
rect 49884 82096 49900 82160
rect 49964 82096 49980 82160
rect 50044 82096 50060 82160
rect 50124 82096 50140 82160
rect 50204 82096 50220 82160
rect 50284 82096 50322 82160
rect 49702 82080 50322 82096
rect 49702 82016 49740 82080
rect 49804 82016 49820 82080
rect 49884 82016 49900 82080
rect 49964 82016 49980 82080
rect 50044 82016 50060 82080
rect 50124 82016 50140 82080
rect 50204 82016 50220 82080
rect 50284 82016 50322 82080
rect 49702 82000 50322 82016
rect 49702 81936 49740 82000
rect 49804 81936 49820 82000
rect 49884 81936 49900 82000
rect 49964 81936 49980 82000
rect 50044 81936 50060 82000
rect 50124 81936 50140 82000
rect 50204 81936 50220 82000
rect 50284 81936 50322 82000
rect 49702 72240 50322 81936
rect 49702 72176 49740 72240
rect 49804 72176 49820 72240
rect 49884 72176 49900 72240
rect 49964 72176 49980 72240
rect 50044 72176 50060 72240
rect 50124 72176 50140 72240
rect 50204 72176 50220 72240
rect 50284 72176 50322 72240
rect 49702 72160 50322 72176
rect 49702 72096 49740 72160
rect 49804 72096 49820 72160
rect 49884 72096 49900 72160
rect 49964 72096 49980 72160
rect 50044 72096 50060 72160
rect 50124 72096 50140 72160
rect 50204 72096 50220 72160
rect 50284 72096 50322 72160
rect 49702 72080 50322 72096
rect 49702 72016 49740 72080
rect 49804 72016 49820 72080
rect 49884 72016 49900 72080
rect 49964 72016 49980 72080
rect 50044 72016 50060 72080
rect 50124 72016 50140 72080
rect 50204 72016 50220 72080
rect 50284 72016 50322 72080
rect 49702 72000 50322 72016
rect 49702 71936 49740 72000
rect 49804 71936 49820 72000
rect 49884 71936 49900 72000
rect 49964 71936 49980 72000
rect 50044 71936 50060 72000
rect 50124 71936 50140 72000
rect 50204 71936 50220 72000
rect 50284 71936 50322 72000
rect 49702 62240 50322 71936
rect 49702 62176 49740 62240
rect 49804 62176 49820 62240
rect 49884 62176 49900 62240
rect 49964 62176 49980 62240
rect 50044 62176 50060 62240
rect 50124 62176 50140 62240
rect 50204 62176 50220 62240
rect 50284 62176 50322 62240
rect 49702 62160 50322 62176
rect 49702 62096 49740 62160
rect 49804 62096 49820 62160
rect 49884 62096 49900 62160
rect 49964 62096 49980 62160
rect 50044 62096 50060 62160
rect 50124 62096 50140 62160
rect 50204 62096 50220 62160
rect 50284 62096 50322 62160
rect 49702 62080 50322 62096
rect 49702 62016 49740 62080
rect 49804 62016 49820 62080
rect 49884 62016 49900 62080
rect 49964 62016 49980 62080
rect 50044 62016 50060 62080
rect 50124 62016 50140 62080
rect 50204 62016 50220 62080
rect 50284 62016 50322 62080
rect 49702 62000 50322 62016
rect 49702 61936 49740 62000
rect 49804 61936 49820 62000
rect 49884 61936 49900 62000
rect 49964 61936 49980 62000
rect 50044 61936 50060 62000
rect 50124 61936 50140 62000
rect 50204 61936 50220 62000
rect 50284 61936 50322 62000
rect 49702 52240 50322 61936
rect 49702 52176 49740 52240
rect 49804 52176 49820 52240
rect 49884 52176 49900 52240
rect 49964 52176 49980 52240
rect 50044 52176 50060 52240
rect 50124 52176 50140 52240
rect 50204 52176 50220 52240
rect 50284 52176 50322 52240
rect 49702 52160 50322 52176
rect 49702 52096 49740 52160
rect 49804 52096 49820 52160
rect 49884 52096 49900 52160
rect 49964 52096 49980 52160
rect 50044 52096 50060 52160
rect 50124 52096 50140 52160
rect 50204 52096 50220 52160
rect 50284 52096 50322 52160
rect 49702 52080 50322 52096
rect 49702 52016 49740 52080
rect 49804 52016 49820 52080
rect 49884 52016 49900 52080
rect 49964 52016 49980 52080
rect 50044 52016 50060 52080
rect 50124 52016 50140 52080
rect 50204 52016 50220 52080
rect 50284 52016 50322 52080
rect 49702 52000 50322 52016
rect 49702 51936 49740 52000
rect 49804 51936 49820 52000
rect 49884 51936 49900 52000
rect 49964 51936 49980 52000
rect 50044 51936 50060 52000
rect 50124 51936 50140 52000
rect 50204 51936 50220 52000
rect 50284 51936 50322 52000
rect 49702 42240 50322 51936
rect 49702 42176 49740 42240
rect 49804 42176 49820 42240
rect 49884 42176 49900 42240
rect 49964 42176 49980 42240
rect 50044 42176 50060 42240
rect 50124 42176 50140 42240
rect 50204 42176 50220 42240
rect 50284 42176 50322 42240
rect 49702 42160 50322 42176
rect 49702 42096 49740 42160
rect 49804 42096 49820 42160
rect 49884 42096 49900 42160
rect 49964 42096 49980 42160
rect 50044 42096 50060 42160
rect 50124 42096 50140 42160
rect 50204 42096 50220 42160
rect 50284 42096 50322 42160
rect 49702 42080 50322 42096
rect 49702 42016 49740 42080
rect 49804 42016 49820 42080
rect 49884 42016 49900 42080
rect 49964 42016 49980 42080
rect 50044 42016 50060 42080
rect 50124 42016 50140 42080
rect 50204 42016 50220 42080
rect 50284 42016 50322 42080
rect 49702 42000 50322 42016
rect 49702 41936 49740 42000
rect 49804 41936 49820 42000
rect 49884 41936 49900 42000
rect 49964 41936 49980 42000
rect 50044 41936 50060 42000
rect 50124 41936 50140 42000
rect 50204 41936 50220 42000
rect 50284 41936 50322 42000
rect 49702 32240 50322 41936
rect 49702 32176 49740 32240
rect 49804 32176 49820 32240
rect 49884 32176 49900 32240
rect 49964 32176 49980 32240
rect 50044 32176 50060 32240
rect 50124 32176 50140 32240
rect 50204 32176 50220 32240
rect 50284 32176 50322 32240
rect 49702 32160 50322 32176
rect 49702 32096 49740 32160
rect 49804 32096 49820 32160
rect 49884 32096 49900 32160
rect 49964 32096 49980 32160
rect 50044 32096 50060 32160
rect 50124 32096 50140 32160
rect 50204 32096 50220 32160
rect 50284 32096 50322 32160
rect 49702 32080 50322 32096
rect 49702 32016 49740 32080
rect 49804 32016 49820 32080
rect 49884 32016 49900 32080
rect 49964 32016 49980 32080
rect 50044 32016 50060 32080
rect 50124 32016 50140 32080
rect 50204 32016 50220 32080
rect 50284 32016 50322 32080
rect 49702 32000 50322 32016
rect 49702 31936 49740 32000
rect 49804 31936 49820 32000
rect 49884 31936 49900 32000
rect 49964 31936 49980 32000
rect 50044 31936 50060 32000
rect 50124 31936 50140 32000
rect 50204 31936 50220 32000
rect 50284 31936 50322 32000
rect 49702 22240 50322 31936
rect 49702 22176 49740 22240
rect 49804 22176 49820 22240
rect 49884 22176 49900 22240
rect 49964 22176 49980 22240
rect 50044 22176 50060 22240
rect 50124 22176 50140 22240
rect 50204 22176 50220 22240
rect 50284 22176 50322 22240
rect 49702 22160 50322 22176
rect 49702 22096 49740 22160
rect 49804 22096 49820 22160
rect 49884 22096 49900 22160
rect 49964 22096 49980 22160
rect 50044 22096 50060 22160
rect 50124 22096 50140 22160
rect 50204 22096 50220 22160
rect 50284 22096 50322 22160
rect 49702 22080 50322 22096
rect 49702 22016 49740 22080
rect 49804 22016 49820 22080
rect 49884 22016 49900 22080
rect 49964 22016 49980 22080
rect 50044 22016 50060 22080
rect 50124 22016 50140 22080
rect 50204 22016 50220 22080
rect 50284 22016 50322 22080
rect 49702 22000 50322 22016
rect 49702 21936 49740 22000
rect 49804 21936 49820 22000
rect 49884 21936 49900 22000
rect 49964 21936 49980 22000
rect 50044 21936 50060 22000
rect 50124 21936 50140 22000
rect 50204 21936 50220 22000
rect 50284 21936 50322 22000
rect 49702 12240 50322 21936
rect 49702 12176 49740 12240
rect 49804 12176 49820 12240
rect 49884 12176 49900 12240
rect 49964 12176 49980 12240
rect 50044 12176 50060 12240
rect 50124 12176 50140 12240
rect 50204 12176 50220 12240
rect 50284 12176 50322 12240
rect 49702 12160 50322 12176
rect 49702 12096 49740 12160
rect 49804 12096 49820 12160
rect 49884 12096 49900 12160
rect 49964 12096 49980 12160
rect 50044 12096 50060 12160
rect 50124 12096 50140 12160
rect 50204 12096 50220 12160
rect 50284 12096 50322 12160
rect 49702 12080 50322 12096
rect 49702 12016 49740 12080
rect 49804 12016 49820 12080
rect 49884 12016 49900 12080
rect 49964 12016 49980 12080
rect 50044 12016 50060 12080
rect 50124 12016 50140 12080
rect 50204 12016 50220 12080
rect 50284 12016 50322 12080
rect 49702 12000 50322 12016
rect 49702 11936 49740 12000
rect 49804 11936 49820 12000
rect 49884 11936 49900 12000
rect 49964 11936 49980 12000
rect 50044 11936 50060 12000
rect 50124 11936 50140 12000
rect 50204 11936 50220 12000
rect 50284 11936 50322 12000
rect 49702 2240 50322 11936
rect 49702 2176 49740 2240
rect 49804 2176 49820 2240
rect 49884 2176 49900 2240
rect 49964 2176 49980 2240
rect 50044 2176 50060 2240
rect 50124 2176 50140 2240
rect 50204 2176 50220 2240
rect 50284 2176 50322 2240
rect 49702 2160 50322 2176
rect 49702 2096 49740 2160
rect 49804 2096 49820 2160
rect 49884 2096 49900 2160
rect 49964 2096 49980 2160
rect 50044 2096 50060 2160
rect 50124 2096 50140 2160
rect 50204 2096 50220 2160
rect 50284 2096 50322 2160
rect 49702 2080 50322 2096
rect 49702 2016 49740 2080
rect 49804 2016 49820 2080
rect 49884 2016 49900 2080
rect 49964 2016 49980 2080
rect 50044 2016 50060 2080
rect 50124 2016 50140 2080
rect 50204 2016 50220 2080
rect 50284 2016 50322 2080
rect 49702 2000 50322 2016
rect 49702 1936 49740 2000
rect 49804 1936 49820 2000
rect 49884 1936 49900 2000
rect 49964 1936 49980 2000
rect 50044 1936 50060 2000
rect 50124 1936 50140 2000
rect 50204 1936 50220 2000
rect 50284 1936 50322 2000
rect 49702 0 50322 1936
rect 52702 84592 53322 87000
rect 52702 84528 52740 84592
rect 52804 84528 52820 84592
rect 52884 84528 52900 84592
rect 52964 84528 52980 84592
rect 53044 84528 53060 84592
rect 53124 84528 53140 84592
rect 53204 84528 53220 84592
rect 53284 84528 53322 84592
rect 52702 84512 53322 84528
rect 52702 84448 52740 84512
rect 52804 84448 52820 84512
rect 52884 84448 52900 84512
rect 52964 84448 52980 84512
rect 53044 84448 53060 84512
rect 53124 84448 53140 84512
rect 53204 84448 53220 84512
rect 53284 84448 53322 84512
rect 52702 84432 53322 84448
rect 52702 84368 52740 84432
rect 52804 84368 52820 84432
rect 52884 84368 52900 84432
rect 52964 84368 52980 84432
rect 53044 84368 53060 84432
rect 53124 84368 53140 84432
rect 53204 84368 53220 84432
rect 53284 84368 53322 84432
rect 52702 84352 53322 84368
rect 52702 84288 52740 84352
rect 52804 84288 52820 84352
rect 52884 84288 52900 84352
rect 52964 84288 52980 84352
rect 53044 84288 53060 84352
rect 53124 84288 53140 84352
rect 53204 84288 53220 84352
rect 53284 84288 53322 84352
rect 52702 74592 53322 84288
rect 52702 74528 52740 74592
rect 52804 74528 52820 74592
rect 52884 74528 52900 74592
rect 52964 74528 52980 74592
rect 53044 74528 53060 74592
rect 53124 74528 53140 74592
rect 53204 74528 53220 74592
rect 53284 74528 53322 74592
rect 52702 74512 53322 74528
rect 52702 74448 52740 74512
rect 52804 74448 52820 74512
rect 52884 74448 52900 74512
rect 52964 74448 52980 74512
rect 53044 74448 53060 74512
rect 53124 74448 53140 74512
rect 53204 74448 53220 74512
rect 53284 74448 53322 74512
rect 52702 74432 53322 74448
rect 52702 74368 52740 74432
rect 52804 74368 52820 74432
rect 52884 74368 52900 74432
rect 52964 74368 52980 74432
rect 53044 74368 53060 74432
rect 53124 74368 53140 74432
rect 53204 74368 53220 74432
rect 53284 74368 53322 74432
rect 52702 74352 53322 74368
rect 52702 74288 52740 74352
rect 52804 74288 52820 74352
rect 52884 74288 52900 74352
rect 52964 74288 52980 74352
rect 53044 74288 53060 74352
rect 53124 74288 53140 74352
rect 53204 74288 53220 74352
rect 53284 74288 53322 74352
rect 52702 64592 53322 74288
rect 52702 64528 52740 64592
rect 52804 64528 52820 64592
rect 52884 64528 52900 64592
rect 52964 64528 52980 64592
rect 53044 64528 53060 64592
rect 53124 64528 53140 64592
rect 53204 64528 53220 64592
rect 53284 64528 53322 64592
rect 52702 64512 53322 64528
rect 52702 64448 52740 64512
rect 52804 64448 52820 64512
rect 52884 64448 52900 64512
rect 52964 64448 52980 64512
rect 53044 64448 53060 64512
rect 53124 64448 53140 64512
rect 53204 64448 53220 64512
rect 53284 64448 53322 64512
rect 52702 64432 53322 64448
rect 52702 64368 52740 64432
rect 52804 64368 52820 64432
rect 52884 64368 52900 64432
rect 52964 64368 52980 64432
rect 53044 64368 53060 64432
rect 53124 64368 53140 64432
rect 53204 64368 53220 64432
rect 53284 64368 53322 64432
rect 52702 64352 53322 64368
rect 52702 64288 52740 64352
rect 52804 64288 52820 64352
rect 52884 64288 52900 64352
rect 52964 64288 52980 64352
rect 53044 64288 53060 64352
rect 53124 64288 53140 64352
rect 53204 64288 53220 64352
rect 53284 64288 53322 64352
rect 52702 54592 53322 64288
rect 52702 54528 52740 54592
rect 52804 54528 52820 54592
rect 52884 54528 52900 54592
rect 52964 54528 52980 54592
rect 53044 54528 53060 54592
rect 53124 54528 53140 54592
rect 53204 54528 53220 54592
rect 53284 54528 53322 54592
rect 52702 54512 53322 54528
rect 52702 54448 52740 54512
rect 52804 54448 52820 54512
rect 52884 54448 52900 54512
rect 52964 54448 52980 54512
rect 53044 54448 53060 54512
rect 53124 54448 53140 54512
rect 53204 54448 53220 54512
rect 53284 54448 53322 54512
rect 52702 54432 53322 54448
rect 52702 54368 52740 54432
rect 52804 54368 52820 54432
rect 52884 54368 52900 54432
rect 52964 54368 52980 54432
rect 53044 54368 53060 54432
rect 53124 54368 53140 54432
rect 53204 54368 53220 54432
rect 53284 54368 53322 54432
rect 52702 54352 53322 54368
rect 52702 54288 52740 54352
rect 52804 54288 52820 54352
rect 52884 54288 52900 54352
rect 52964 54288 52980 54352
rect 53044 54288 53060 54352
rect 53124 54288 53140 54352
rect 53204 54288 53220 54352
rect 53284 54288 53322 54352
rect 52702 44592 53322 54288
rect 52702 44528 52740 44592
rect 52804 44528 52820 44592
rect 52884 44528 52900 44592
rect 52964 44528 52980 44592
rect 53044 44528 53060 44592
rect 53124 44528 53140 44592
rect 53204 44528 53220 44592
rect 53284 44528 53322 44592
rect 52702 44512 53322 44528
rect 52702 44448 52740 44512
rect 52804 44448 52820 44512
rect 52884 44448 52900 44512
rect 52964 44448 52980 44512
rect 53044 44448 53060 44512
rect 53124 44448 53140 44512
rect 53204 44448 53220 44512
rect 53284 44448 53322 44512
rect 52702 44432 53322 44448
rect 52702 44368 52740 44432
rect 52804 44368 52820 44432
rect 52884 44368 52900 44432
rect 52964 44368 52980 44432
rect 53044 44368 53060 44432
rect 53124 44368 53140 44432
rect 53204 44368 53220 44432
rect 53284 44368 53322 44432
rect 52702 44352 53322 44368
rect 52702 44288 52740 44352
rect 52804 44288 52820 44352
rect 52884 44288 52900 44352
rect 52964 44288 52980 44352
rect 53044 44288 53060 44352
rect 53124 44288 53140 44352
rect 53204 44288 53220 44352
rect 53284 44288 53322 44352
rect 52702 34592 53322 44288
rect 52702 34528 52740 34592
rect 52804 34528 52820 34592
rect 52884 34528 52900 34592
rect 52964 34528 52980 34592
rect 53044 34528 53060 34592
rect 53124 34528 53140 34592
rect 53204 34528 53220 34592
rect 53284 34528 53322 34592
rect 52702 34512 53322 34528
rect 52702 34448 52740 34512
rect 52804 34448 52820 34512
rect 52884 34448 52900 34512
rect 52964 34448 52980 34512
rect 53044 34448 53060 34512
rect 53124 34448 53140 34512
rect 53204 34448 53220 34512
rect 53284 34448 53322 34512
rect 52702 34432 53322 34448
rect 52702 34368 52740 34432
rect 52804 34368 52820 34432
rect 52884 34368 52900 34432
rect 52964 34368 52980 34432
rect 53044 34368 53060 34432
rect 53124 34368 53140 34432
rect 53204 34368 53220 34432
rect 53284 34368 53322 34432
rect 52702 34352 53322 34368
rect 52702 34288 52740 34352
rect 52804 34288 52820 34352
rect 52884 34288 52900 34352
rect 52964 34288 52980 34352
rect 53044 34288 53060 34352
rect 53124 34288 53140 34352
rect 53204 34288 53220 34352
rect 53284 34288 53322 34352
rect 52702 24592 53322 34288
rect 52702 24528 52740 24592
rect 52804 24528 52820 24592
rect 52884 24528 52900 24592
rect 52964 24528 52980 24592
rect 53044 24528 53060 24592
rect 53124 24528 53140 24592
rect 53204 24528 53220 24592
rect 53284 24528 53322 24592
rect 52702 24512 53322 24528
rect 52702 24448 52740 24512
rect 52804 24448 52820 24512
rect 52884 24448 52900 24512
rect 52964 24448 52980 24512
rect 53044 24448 53060 24512
rect 53124 24448 53140 24512
rect 53204 24448 53220 24512
rect 53284 24448 53322 24512
rect 52702 24432 53322 24448
rect 52702 24368 52740 24432
rect 52804 24368 52820 24432
rect 52884 24368 52900 24432
rect 52964 24368 52980 24432
rect 53044 24368 53060 24432
rect 53124 24368 53140 24432
rect 53204 24368 53220 24432
rect 53284 24368 53322 24432
rect 52702 24352 53322 24368
rect 52702 24288 52740 24352
rect 52804 24288 52820 24352
rect 52884 24288 52900 24352
rect 52964 24288 52980 24352
rect 53044 24288 53060 24352
rect 53124 24288 53140 24352
rect 53204 24288 53220 24352
rect 53284 24288 53322 24352
rect 52702 14592 53322 24288
rect 52702 14528 52740 14592
rect 52804 14528 52820 14592
rect 52884 14528 52900 14592
rect 52964 14528 52980 14592
rect 53044 14528 53060 14592
rect 53124 14528 53140 14592
rect 53204 14528 53220 14592
rect 53284 14528 53322 14592
rect 52702 14512 53322 14528
rect 52702 14448 52740 14512
rect 52804 14448 52820 14512
rect 52884 14448 52900 14512
rect 52964 14448 52980 14512
rect 53044 14448 53060 14512
rect 53124 14448 53140 14512
rect 53204 14448 53220 14512
rect 53284 14448 53322 14512
rect 52702 14432 53322 14448
rect 52702 14368 52740 14432
rect 52804 14368 52820 14432
rect 52884 14368 52900 14432
rect 52964 14368 52980 14432
rect 53044 14368 53060 14432
rect 53124 14368 53140 14432
rect 53204 14368 53220 14432
rect 53284 14368 53322 14432
rect 52702 14352 53322 14368
rect 52702 14288 52740 14352
rect 52804 14288 52820 14352
rect 52884 14288 52900 14352
rect 52964 14288 52980 14352
rect 53044 14288 53060 14352
rect 53124 14288 53140 14352
rect 53204 14288 53220 14352
rect 53284 14288 53322 14352
rect 52702 4592 53322 14288
rect 52702 4528 52740 4592
rect 52804 4528 52820 4592
rect 52884 4528 52900 4592
rect 52964 4528 52980 4592
rect 53044 4528 53060 4592
rect 53124 4528 53140 4592
rect 53204 4528 53220 4592
rect 53284 4528 53322 4592
rect 52702 4512 53322 4528
rect 52702 4448 52740 4512
rect 52804 4448 52820 4512
rect 52884 4448 52900 4512
rect 52964 4448 52980 4512
rect 53044 4448 53060 4512
rect 53124 4448 53140 4512
rect 53204 4448 53220 4512
rect 53284 4448 53322 4512
rect 52702 4432 53322 4448
rect 52702 4368 52740 4432
rect 52804 4368 52820 4432
rect 52884 4368 52900 4432
rect 52964 4368 52980 4432
rect 53044 4368 53060 4432
rect 53124 4368 53140 4432
rect 53204 4368 53220 4432
rect 53284 4368 53322 4432
rect 52702 4352 53322 4368
rect 52702 4288 52740 4352
rect 52804 4288 52820 4352
rect 52884 4288 52900 4352
rect 52964 4288 52980 4352
rect 53044 4288 53060 4352
rect 53124 4288 53140 4352
rect 53204 4288 53220 4352
rect 53284 4288 53322 4352
rect 52702 0 53322 4288
rect 55702 82240 56322 87000
rect 55702 82176 55740 82240
rect 55804 82176 55820 82240
rect 55884 82176 55900 82240
rect 55964 82176 55980 82240
rect 56044 82176 56060 82240
rect 56124 82176 56140 82240
rect 56204 82176 56220 82240
rect 56284 82176 56322 82240
rect 55702 82160 56322 82176
rect 55702 82096 55740 82160
rect 55804 82096 55820 82160
rect 55884 82096 55900 82160
rect 55964 82096 55980 82160
rect 56044 82096 56060 82160
rect 56124 82096 56140 82160
rect 56204 82096 56220 82160
rect 56284 82096 56322 82160
rect 55702 82080 56322 82096
rect 55702 82016 55740 82080
rect 55804 82016 55820 82080
rect 55884 82016 55900 82080
rect 55964 82016 55980 82080
rect 56044 82016 56060 82080
rect 56124 82016 56140 82080
rect 56204 82016 56220 82080
rect 56284 82016 56322 82080
rect 55702 82000 56322 82016
rect 55702 81936 55740 82000
rect 55804 81936 55820 82000
rect 55884 81936 55900 82000
rect 55964 81936 55980 82000
rect 56044 81936 56060 82000
rect 56124 81936 56140 82000
rect 56204 81936 56220 82000
rect 56284 81936 56322 82000
rect 55702 72240 56322 81936
rect 55702 72176 55740 72240
rect 55804 72176 55820 72240
rect 55884 72176 55900 72240
rect 55964 72176 55980 72240
rect 56044 72176 56060 72240
rect 56124 72176 56140 72240
rect 56204 72176 56220 72240
rect 56284 72176 56322 72240
rect 55702 72160 56322 72176
rect 55702 72096 55740 72160
rect 55804 72096 55820 72160
rect 55884 72096 55900 72160
rect 55964 72096 55980 72160
rect 56044 72096 56060 72160
rect 56124 72096 56140 72160
rect 56204 72096 56220 72160
rect 56284 72096 56322 72160
rect 55702 72080 56322 72096
rect 55702 72016 55740 72080
rect 55804 72016 55820 72080
rect 55884 72016 55900 72080
rect 55964 72016 55980 72080
rect 56044 72016 56060 72080
rect 56124 72016 56140 72080
rect 56204 72016 56220 72080
rect 56284 72016 56322 72080
rect 55702 72000 56322 72016
rect 55702 71936 55740 72000
rect 55804 71936 55820 72000
rect 55884 71936 55900 72000
rect 55964 71936 55980 72000
rect 56044 71936 56060 72000
rect 56124 71936 56140 72000
rect 56204 71936 56220 72000
rect 56284 71936 56322 72000
rect 55702 62240 56322 71936
rect 55702 62176 55740 62240
rect 55804 62176 55820 62240
rect 55884 62176 55900 62240
rect 55964 62176 55980 62240
rect 56044 62176 56060 62240
rect 56124 62176 56140 62240
rect 56204 62176 56220 62240
rect 56284 62176 56322 62240
rect 55702 62160 56322 62176
rect 55702 62096 55740 62160
rect 55804 62096 55820 62160
rect 55884 62096 55900 62160
rect 55964 62096 55980 62160
rect 56044 62096 56060 62160
rect 56124 62096 56140 62160
rect 56204 62096 56220 62160
rect 56284 62096 56322 62160
rect 55702 62080 56322 62096
rect 55702 62016 55740 62080
rect 55804 62016 55820 62080
rect 55884 62016 55900 62080
rect 55964 62016 55980 62080
rect 56044 62016 56060 62080
rect 56124 62016 56140 62080
rect 56204 62016 56220 62080
rect 56284 62016 56322 62080
rect 55702 62000 56322 62016
rect 55702 61936 55740 62000
rect 55804 61936 55820 62000
rect 55884 61936 55900 62000
rect 55964 61936 55980 62000
rect 56044 61936 56060 62000
rect 56124 61936 56140 62000
rect 56204 61936 56220 62000
rect 56284 61936 56322 62000
rect 55702 52240 56322 61936
rect 55702 52176 55740 52240
rect 55804 52176 55820 52240
rect 55884 52176 55900 52240
rect 55964 52176 55980 52240
rect 56044 52176 56060 52240
rect 56124 52176 56140 52240
rect 56204 52176 56220 52240
rect 56284 52176 56322 52240
rect 55702 52160 56322 52176
rect 55702 52096 55740 52160
rect 55804 52096 55820 52160
rect 55884 52096 55900 52160
rect 55964 52096 55980 52160
rect 56044 52096 56060 52160
rect 56124 52096 56140 52160
rect 56204 52096 56220 52160
rect 56284 52096 56322 52160
rect 55702 52080 56322 52096
rect 55702 52016 55740 52080
rect 55804 52016 55820 52080
rect 55884 52016 55900 52080
rect 55964 52016 55980 52080
rect 56044 52016 56060 52080
rect 56124 52016 56140 52080
rect 56204 52016 56220 52080
rect 56284 52016 56322 52080
rect 55702 52000 56322 52016
rect 55702 51936 55740 52000
rect 55804 51936 55820 52000
rect 55884 51936 55900 52000
rect 55964 51936 55980 52000
rect 56044 51936 56060 52000
rect 56124 51936 56140 52000
rect 56204 51936 56220 52000
rect 56284 51936 56322 52000
rect 55702 42240 56322 51936
rect 55702 42176 55740 42240
rect 55804 42176 55820 42240
rect 55884 42176 55900 42240
rect 55964 42176 55980 42240
rect 56044 42176 56060 42240
rect 56124 42176 56140 42240
rect 56204 42176 56220 42240
rect 56284 42176 56322 42240
rect 55702 42160 56322 42176
rect 55702 42096 55740 42160
rect 55804 42096 55820 42160
rect 55884 42096 55900 42160
rect 55964 42096 55980 42160
rect 56044 42096 56060 42160
rect 56124 42096 56140 42160
rect 56204 42096 56220 42160
rect 56284 42096 56322 42160
rect 55702 42080 56322 42096
rect 55702 42016 55740 42080
rect 55804 42016 55820 42080
rect 55884 42016 55900 42080
rect 55964 42016 55980 42080
rect 56044 42016 56060 42080
rect 56124 42016 56140 42080
rect 56204 42016 56220 42080
rect 56284 42016 56322 42080
rect 55702 42000 56322 42016
rect 55702 41936 55740 42000
rect 55804 41936 55820 42000
rect 55884 41936 55900 42000
rect 55964 41936 55980 42000
rect 56044 41936 56060 42000
rect 56124 41936 56140 42000
rect 56204 41936 56220 42000
rect 56284 41936 56322 42000
rect 55702 32240 56322 41936
rect 55702 32176 55740 32240
rect 55804 32176 55820 32240
rect 55884 32176 55900 32240
rect 55964 32176 55980 32240
rect 56044 32176 56060 32240
rect 56124 32176 56140 32240
rect 56204 32176 56220 32240
rect 56284 32176 56322 32240
rect 55702 32160 56322 32176
rect 55702 32096 55740 32160
rect 55804 32096 55820 32160
rect 55884 32096 55900 32160
rect 55964 32096 55980 32160
rect 56044 32096 56060 32160
rect 56124 32096 56140 32160
rect 56204 32096 56220 32160
rect 56284 32096 56322 32160
rect 55702 32080 56322 32096
rect 55702 32016 55740 32080
rect 55804 32016 55820 32080
rect 55884 32016 55900 32080
rect 55964 32016 55980 32080
rect 56044 32016 56060 32080
rect 56124 32016 56140 32080
rect 56204 32016 56220 32080
rect 56284 32016 56322 32080
rect 55702 32000 56322 32016
rect 55702 31936 55740 32000
rect 55804 31936 55820 32000
rect 55884 31936 55900 32000
rect 55964 31936 55980 32000
rect 56044 31936 56060 32000
rect 56124 31936 56140 32000
rect 56204 31936 56220 32000
rect 56284 31936 56322 32000
rect 55702 22240 56322 31936
rect 55702 22176 55740 22240
rect 55804 22176 55820 22240
rect 55884 22176 55900 22240
rect 55964 22176 55980 22240
rect 56044 22176 56060 22240
rect 56124 22176 56140 22240
rect 56204 22176 56220 22240
rect 56284 22176 56322 22240
rect 55702 22160 56322 22176
rect 55702 22096 55740 22160
rect 55804 22096 55820 22160
rect 55884 22096 55900 22160
rect 55964 22096 55980 22160
rect 56044 22096 56060 22160
rect 56124 22096 56140 22160
rect 56204 22096 56220 22160
rect 56284 22096 56322 22160
rect 55702 22080 56322 22096
rect 55702 22016 55740 22080
rect 55804 22016 55820 22080
rect 55884 22016 55900 22080
rect 55964 22016 55980 22080
rect 56044 22016 56060 22080
rect 56124 22016 56140 22080
rect 56204 22016 56220 22080
rect 56284 22016 56322 22080
rect 55702 22000 56322 22016
rect 55702 21936 55740 22000
rect 55804 21936 55820 22000
rect 55884 21936 55900 22000
rect 55964 21936 55980 22000
rect 56044 21936 56060 22000
rect 56124 21936 56140 22000
rect 56204 21936 56220 22000
rect 56284 21936 56322 22000
rect 55702 12240 56322 21936
rect 55702 12176 55740 12240
rect 55804 12176 55820 12240
rect 55884 12176 55900 12240
rect 55964 12176 55980 12240
rect 56044 12176 56060 12240
rect 56124 12176 56140 12240
rect 56204 12176 56220 12240
rect 56284 12176 56322 12240
rect 55702 12160 56322 12176
rect 55702 12096 55740 12160
rect 55804 12096 55820 12160
rect 55884 12096 55900 12160
rect 55964 12096 55980 12160
rect 56044 12096 56060 12160
rect 56124 12096 56140 12160
rect 56204 12096 56220 12160
rect 56284 12096 56322 12160
rect 55702 12080 56322 12096
rect 55702 12016 55740 12080
rect 55804 12016 55820 12080
rect 55884 12016 55900 12080
rect 55964 12016 55980 12080
rect 56044 12016 56060 12080
rect 56124 12016 56140 12080
rect 56204 12016 56220 12080
rect 56284 12016 56322 12080
rect 55702 12000 56322 12016
rect 55702 11936 55740 12000
rect 55804 11936 55820 12000
rect 55884 11936 55900 12000
rect 55964 11936 55980 12000
rect 56044 11936 56060 12000
rect 56124 11936 56140 12000
rect 56204 11936 56220 12000
rect 56284 11936 56322 12000
rect 55702 2240 56322 11936
rect 55702 2176 55740 2240
rect 55804 2176 55820 2240
rect 55884 2176 55900 2240
rect 55964 2176 55980 2240
rect 56044 2176 56060 2240
rect 56124 2176 56140 2240
rect 56204 2176 56220 2240
rect 56284 2176 56322 2240
rect 55702 2160 56322 2176
rect 55702 2096 55740 2160
rect 55804 2096 55820 2160
rect 55884 2096 55900 2160
rect 55964 2096 55980 2160
rect 56044 2096 56060 2160
rect 56124 2096 56140 2160
rect 56204 2096 56220 2160
rect 56284 2096 56322 2160
rect 55702 2080 56322 2096
rect 55702 2016 55740 2080
rect 55804 2016 55820 2080
rect 55884 2016 55900 2080
rect 55964 2016 55980 2080
rect 56044 2016 56060 2080
rect 56124 2016 56140 2080
rect 56204 2016 56220 2080
rect 56284 2016 56322 2080
rect 55702 2000 56322 2016
rect 55702 1936 55740 2000
rect 55804 1936 55820 2000
rect 55884 1936 55900 2000
rect 55964 1936 55980 2000
rect 56044 1936 56060 2000
rect 56124 1936 56140 2000
rect 56204 1936 56220 2000
rect 56284 1936 56322 2000
rect 55702 0 56322 1936
rect 58702 84592 59322 87000
rect 58702 84528 58740 84592
rect 58804 84528 58820 84592
rect 58884 84528 58900 84592
rect 58964 84528 58980 84592
rect 59044 84528 59060 84592
rect 59124 84528 59140 84592
rect 59204 84528 59220 84592
rect 59284 84528 59322 84592
rect 58702 84512 59322 84528
rect 58702 84448 58740 84512
rect 58804 84448 58820 84512
rect 58884 84448 58900 84512
rect 58964 84448 58980 84512
rect 59044 84448 59060 84512
rect 59124 84448 59140 84512
rect 59204 84448 59220 84512
rect 59284 84448 59322 84512
rect 58702 84432 59322 84448
rect 58702 84368 58740 84432
rect 58804 84368 58820 84432
rect 58884 84368 58900 84432
rect 58964 84368 58980 84432
rect 59044 84368 59060 84432
rect 59124 84368 59140 84432
rect 59204 84368 59220 84432
rect 59284 84368 59322 84432
rect 58702 84352 59322 84368
rect 58702 84288 58740 84352
rect 58804 84288 58820 84352
rect 58884 84288 58900 84352
rect 58964 84288 58980 84352
rect 59044 84288 59060 84352
rect 59124 84288 59140 84352
rect 59204 84288 59220 84352
rect 59284 84288 59322 84352
rect 58702 74592 59322 84288
rect 58702 74528 58740 74592
rect 58804 74528 58820 74592
rect 58884 74528 58900 74592
rect 58964 74528 58980 74592
rect 59044 74528 59060 74592
rect 59124 74528 59140 74592
rect 59204 74528 59220 74592
rect 59284 74528 59322 74592
rect 58702 74512 59322 74528
rect 58702 74448 58740 74512
rect 58804 74448 58820 74512
rect 58884 74448 58900 74512
rect 58964 74448 58980 74512
rect 59044 74448 59060 74512
rect 59124 74448 59140 74512
rect 59204 74448 59220 74512
rect 59284 74448 59322 74512
rect 58702 74432 59322 74448
rect 58702 74368 58740 74432
rect 58804 74368 58820 74432
rect 58884 74368 58900 74432
rect 58964 74368 58980 74432
rect 59044 74368 59060 74432
rect 59124 74368 59140 74432
rect 59204 74368 59220 74432
rect 59284 74368 59322 74432
rect 58702 74352 59322 74368
rect 58702 74288 58740 74352
rect 58804 74288 58820 74352
rect 58884 74288 58900 74352
rect 58964 74288 58980 74352
rect 59044 74288 59060 74352
rect 59124 74288 59140 74352
rect 59204 74288 59220 74352
rect 59284 74288 59322 74352
rect 58702 64592 59322 74288
rect 58702 64528 58740 64592
rect 58804 64528 58820 64592
rect 58884 64528 58900 64592
rect 58964 64528 58980 64592
rect 59044 64528 59060 64592
rect 59124 64528 59140 64592
rect 59204 64528 59220 64592
rect 59284 64528 59322 64592
rect 58702 64512 59322 64528
rect 58702 64448 58740 64512
rect 58804 64448 58820 64512
rect 58884 64448 58900 64512
rect 58964 64448 58980 64512
rect 59044 64448 59060 64512
rect 59124 64448 59140 64512
rect 59204 64448 59220 64512
rect 59284 64448 59322 64512
rect 58702 64432 59322 64448
rect 58702 64368 58740 64432
rect 58804 64368 58820 64432
rect 58884 64368 58900 64432
rect 58964 64368 58980 64432
rect 59044 64368 59060 64432
rect 59124 64368 59140 64432
rect 59204 64368 59220 64432
rect 59284 64368 59322 64432
rect 58702 64352 59322 64368
rect 58702 64288 58740 64352
rect 58804 64288 58820 64352
rect 58884 64288 58900 64352
rect 58964 64288 58980 64352
rect 59044 64288 59060 64352
rect 59124 64288 59140 64352
rect 59204 64288 59220 64352
rect 59284 64288 59322 64352
rect 58702 54592 59322 64288
rect 58702 54528 58740 54592
rect 58804 54528 58820 54592
rect 58884 54528 58900 54592
rect 58964 54528 58980 54592
rect 59044 54528 59060 54592
rect 59124 54528 59140 54592
rect 59204 54528 59220 54592
rect 59284 54528 59322 54592
rect 58702 54512 59322 54528
rect 58702 54448 58740 54512
rect 58804 54448 58820 54512
rect 58884 54448 58900 54512
rect 58964 54448 58980 54512
rect 59044 54448 59060 54512
rect 59124 54448 59140 54512
rect 59204 54448 59220 54512
rect 59284 54448 59322 54512
rect 58702 54432 59322 54448
rect 58702 54368 58740 54432
rect 58804 54368 58820 54432
rect 58884 54368 58900 54432
rect 58964 54368 58980 54432
rect 59044 54368 59060 54432
rect 59124 54368 59140 54432
rect 59204 54368 59220 54432
rect 59284 54368 59322 54432
rect 58702 54352 59322 54368
rect 58702 54288 58740 54352
rect 58804 54288 58820 54352
rect 58884 54288 58900 54352
rect 58964 54288 58980 54352
rect 59044 54288 59060 54352
rect 59124 54288 59140 54352
rect 59204 54288 59220 54352
rect 59284 54288 59322 54352
rect 58702 44592 59322 54288
rect 58702 44528 58740 44592
rect 58804 44528 58820 44592
rect 58884 44528 58900 44592
rect 58964 44528 58980 44592
rect 59044 44528 59060 44592
rect 59124 44528 59140 44592
rect 59204 44528 59220 44592
rect 59284 44528 59322 44592
rect 58702 44512 59322 44528
rect 58702 44448 58740 44512
rect 58804 44448 58820 44512
rect 58884 44448 58900 44512
rect 58964 44448 58980 44512
rect 59044 44448 59060 44512
rect 59124 44448 59140 44512
rect 59204 44448 59220 44512
rect 59284 44448 59322 44512
rect 58702 44432 59322 44448
rect 58702 44368 58740 44432
rect 58804 44368 58820 44432
rect 58884 44368 58900 44432
rect 58964 44368 58980 44432
rect 59044 44368 59060 44432
rect 59124 44368 59140 44432
rect 59204 44368 59220 44432
rect 59284 44368 59322 44432
rect 58702 44352 59322 44368
rect 58702 44288 58740 44352
rect 58804 44288 58820 44352
rect 58884 44288 58900 44352
rect 58964 44288 58980 44352
rect 59044 44288 59060 44352
rect 59124 44288 59140 44352
rect 59204 44288 59220 44352
rect 59284 44288 59322 44352
rect 58702 34592 59322 44288
rect 58702 34528 58740 34592
rect 58804 34528 58820 34592
rect 58884 34528 58900 34592
rect 58964 34528 58980 34592
rect 59044 34528 59060 34592
rect 59124 34528 59140 34592
rect 59204 34528 59220 34592
rect 59284 34528 59322 34592
rect 58702 34512 59322 34528
rect 58702 34448 58740 34512
rect 58804 34448 58820 34512
rect 58884 34448 58900 34512
rect 58964 34448 58980 34512
rect 59044 34448 59060 34512
rect 59124 34448 59140 34512
rect 59204 34448 59220 34512
rect 59284 34448 59322 34512
rect 58702 34432 59322 34448
rect 58702 34368 58740 34432
rect 58804 34368 58820 34432
rect 58884 34368 58900 34432
rect 58964 34368 58980 34432
rect 59044 34368 59060 34432
rect 59124 34368 59140 34432
rect 59204 34368 59220 34432
rect 59284 34368 59322 34432
rect 58702 34352 59322 34368
rect 58702 34288 58740 34352
rect 58804 34288 58820 34352
rect 58884 34288 58900 34352
rect 58964 34288 58980 34352
rect 59044 34288 59060 34352
rect 59124 34288 59140 34352
rect 59204 34288 59220 34352
rect 59284 34288 59322 34352
rect 58702 24592 59322 34288
rect 58702 24528 58740 24592
rect 58804 24528 58820 24592
rect 58884 24528 58900 24592
rect 58964 24528 58980 24592
rect 59044 24528 59060 24592
rect 59124 24528 59140 24592
rect 59204 24528 59220 24592
rect 59284 24528 59322 24592
rect 58702 24512 59322 24528
rect 58702 24448 58740 24512
rect 58804 24448 58820 24512
rect 58884 24448 58900 24512
rect 58964 24448 58980 24512
rect 59044 24448 59060 24512
rect 59124 24448 59140 24512
rect 59204 24448 59220 24512
rect 59284 24448 59322 24512
rect 58702 24432 59322 24448
rect 58702 24368 58740 24432
rect 58804 24368 58820 24432
rect 58884 24368 58900 24432
rect 58964 24368 58980 24432
rect 59044 24368 59060 24432
rect 59124 24368 59140 24432
rect 59204 24368 59220 24432
rect 59284 24368 59322 24432
rect 58702 24352 59322 24368
rect 58702 24288 58740 24352
rect 58804 24288 58820 24352
rect 58884 24288 58900 24352
rect 58964 24288 58980 24352
rect 59044 24288 59060 24352
rect 59124 24288 59140 24352
rect 59204 24288 59220 24352
rect 59284 24288 59322 24352
rect 58702 14592 59322 24288
rect 58702 14528 58740 14592
rect 58804 14528 58820 14592
rect 58884 14528 58900 14592
rect 58964 14528 58980 14592
rect 59044 14528 59060 14592
rect 59124 14528 59140 14592
rect 59204 14528 59220 14592
rect 59284 14528 59322 14592
rect 58702 14512 59322 14528
rect 58702 14448 58740 14512
rect 58804 14448 58820 14512
rect 58884 14448 58900 14512
rect 58964 14448 58980 14512
rect 59044 14448 59060 14512
rect 59124 14448 59140 14512
rect 59204 14448 59220 14512
rect 59284 14448 59322 14512
rect 58702 14432 59322 14448
rect 58702 14368 58740 14432
rect 58804 14368 58820 14432
rect 58884 14368 58900 14432
rect 58964 14368 58980 14432
rect 59044 14368 59060 14432
rect 59124 14368 59140 14432
rect 59204 14368 59220 14432
rect 59284 14368 59322 14432
rect 58702 14352 59322 14368
rect 58702 14288 58740 14352
rect 58804 14288 58820 14352
rect 58884 14288 58900 14352
rect 58964 14288 58980 14352
rect 59044 14288 59060 14352
rect 59124 14288 59140 14352
rect 59204 14288 59220 14352
rect 59284 14288 59322 14352
rect 58702 4592 59322 14288
rect 58702 4528 58740 4592
rect 58804 4528 58820 4592
rect 58884 4528 58900 4592
rect 58964 4528 58980 4592
rect 59044 4528 59060 4592
rect 59124 4528 59140 4592
rect 59204 4528 59220 4592
rect 59284 4528 59322 4592
rect 58702 4512 59322 4528
rect 58702 4448 58740 4512
rect 58804 4448 58820 4512
rect 58884 4448 58900 4512
rect 58964 4448 58980 4512
rect 59044 4448 59060 4512
rect 59124 4448 59140 4512
rect 59204 4448 59220 4512
rect 59284 4448 59322 4512
rect 58702 4432 59322 4448
rect 58702 4368 58740 4432
rect 58804 4368 58820 4432
rect 58884 4368 58900 4432
rect 58964 4368 58980 4432
rect 59044 4368 59060 4432
rect 59124 4368 59140 4432
rect 59204 4368 59220 4432
rect 59284 4368 59322 4432
rect 58702 4352 59322 4368
rect 58702 4288 58740 4352
rect 58804 4288 58820 4352
rect 58884 4288 58900 4352
rect 58964 4288 58980 4352
rect 59044 4288 59060 4352
rect 59124 4288 59140 4352
rect 59204 4288 59220 4352
rect 59284 4288 59322 4352
rect 58702 0 59322 4288
rect 61702 82240 62322 87000
rect 61702 82176 61740 82240
rect 61804 82176 61820 82240
rect 61884 82176 61900 82240
rect 61964 82176 61980 82240
rect 62044 82176 62060 82240
rect 62124 82176 62140 82240
rect 62204 82176 62220 82240
rect 62284 82176 62322 82240
rect 61702 82160 62322 82176
rect 61702 82096 61740 82160
rect 61804 82096 61820 82160
rect 61884 82096 61900 82160
rect 61964 82096 61980 82160
rect 62044 82096 62060 82160
rect 62124 82096 62140 82160
rect 62204 82096 62220 82160
rect 62284 82096 62322 82160
rect 61702 82080 62322 82096
rect 61702 82016 61740 82080
rect 61804 82016 61820 82080
rect 61884 82016 61900 82080
rect 61964 82016 61980 82080
rect 62044 82016 62060 82080
rect 62124 82016 62140 82080
rect 62204 82016 62220 82080
rect 62284 82016 62322 82080
rect 61702 82000 62322 82016
rect 61702 81936 61740 82000
rect 61804 81936 61820 82000
rect 61884 81936 61900 82000
rect 61964 81936 61980 82000
rect 62044 81936 62060 82000
rect 62124 81936 62140 82000
rect 62204 81936 62220 82000
rect 62284 81936 62322 82000
rect 61702 72240 62322 81936
rect 61702 72176 61740 72240
rect 61804 72176 61820 72240
rect 61884 72176 61900 72240
rect 61964 72176 61980 72240
rect 62044 72176 62060 72240
rect 62124 72176 62140 72240
rect 62204 72176 62220 72240
rect 62284 72176 62322 72240
rect 61702 72160 62322 72176
rect 61702 72096 61740 72160
rect 61804 72096 61820 72160
rect 61884 72096 61900 72160
rect 61964 72096 61980 72160
rect 62044 72096 62060 72160
rect 62124 72096 62140 72160
rect 62204 72096 62220 72160
rect 62284 72096 62322 72160
rect 61702 72080 62322 72096
rect 61702 72016 61740 72080
rect 61804 72016 61820 72080
rect 61884 72016 61900 72080
rect 61964 72016 61980 72080
rect 62044 72016 62060 72080
rect 62124 72016 62140 72080
rect 62204 72016 62220 72080
rect 62284 72016 62322 72080
rect 61702 72000 62322 72016
rect 61702 71936 61740 72000
rect 61804 71936 61820 72000
rect 61884 71936 61900 72000
rect 61964 71936 61980 72000
rect 62044 71936 62060 72000
rect 62124 71936 62140 72000
rect 62204 71936 62220 72000
rect 62284 71936 62322 72000
rect 61702 62240 62322 71936
rect 64702 84592 65322 87000
rect 64702 84528 64740 84592
rect 64804 84528 64820 84592
rect 64884 84528 64900 84592
rect 64964 84528 64980 84592
rect 65044 84528 65060 84592
rect 65124 84528 65140 84592
rect 65204 84528 65220 84592
rect 65284 84528 65322 84592
rect 64702 84512 65322 84528
rect 64702 84448 64740 84512
rect 64804 84448 64820 84512
rect 64884 84448 64900 84512
rect 64964 84448 64980 84512
rect 65044 84448 65060 84512
rect 65124 84448 65140 84512
rect 65204 84448 65220 84512
rect 65284 84448 65322 84512
rect 64702 84432 65322 84448
rect 64702 84368 64740 84432
rect 64804 84368 64820 84432
rect 64884 84368 64900 84432
rect 64964 84368 64980 84432
rect 65044 84368 65060 84432
rect 65124 84368 65140 84432
rect 65204 84368 65220 84432
rect 65284 84368 65322 84432
rect 64702 84352 65322 84368
rect 64702 84288 64740 84352
rect 64804 84288 64820 84352
rect 64884 84288 64900 84352
rect 64964 84288 64980 84352
rect 65044 84288 65060 84352
rect 65124 84288 65140 84352
rect 65204 84288 65220 84352
rect 65284 84288 65322 84352
rect 64702 74592 65322 84288
rect 64702 74528 64740 74592
rect 64804 74528 64820 74592
rect 64884 74528 64900 74592
rect 64964 74528 64980 74592
rect 65044 74528 65060 74592
rect 65124 74528 65140 74592
rect 65204 74528 65220 74592
rect 65284 74528 65322 74592
rect 64702 74512 65322 74528
rect 64702 74448 64740 74512
rect 64804 74448 64820 74512
rect 64884 74448 64900 74512
rect 64964 74448 64980 74512
rect 65044 74448 65060 74512
rect 65124 74448 65140 74512
rect 65204 74448 65220 74512
rect 65284 74448 65322 74512
rect 64702 74432 65322 74448
rect 64702 74368 64740 74432
rect 64804 74368 64820 74432
rect 64884 74368 64900 74432
rect 64964 74368 64980 74432
rect 65044 74368 65060 74432
rect 65124 74368 65140 74432
rect 65204 74368 65220 74432
rect 65284 74368 65322 74432
rect 64702 74352 65322 74368
rect 64702 74288 64740 74352
rect 64804 74288 64820 74352
rect 64884 74288 64900 74352
rect 64964 74288 64980 74352
rect 65044 74288 65060 74352
rect 65124 74288 65140 74352
rect 65204 74288 65220 74352
rect 65284 74288 65322 74352
rect 63539 65244 63605 65245
rect 63539 65180 63540 65244
rect 63604 65180 63605 65244
rect 63539 65179 63605 65180
rect 61702 62176 61740 62240
rect 61804 62176 61820 62240
rect 61884 62176 61900 62240
rect 61964 62176 61980 62240
rect 62044 62176 62060 62240
rect 62124 62176 62140 62240
rect 62204 62176 62220 62240
rect 62284 62176 62322 62240
rect 61702 62160 62322 62176
rect 61702 62096 61740 62160
rect 61804 62096 61820 62160
rect 61884 62096 61900 62160
rect 61964 62096 61980 62160
rect 62044 62096 62060 62160
rect 62124 62096 62140 62160
rect 62204 62096 62220 62160
rect 62284 62096 62322 62160
rect 61702 62080 62322 62096
rect 61702 62016 61740 62080
rect 61804 62016 61820 62080
rect 61884 62016 61900 62080
rect 61964 62016 61980 62080
rect 62044 62016 62060 62080
rect 62124 62016 62140 62080
rect 62204 62016 62220 62080
rect 62284 62016 62322 62080
rect 61702 62000 62322 62016
rect 61702 61936 61740 62000
rect 61804 61936 61820 62000
rect 61884 61936 61900 62000
rect 61964 61936 61980 62000
rect 62044 61936 62060 62000
rect 62124 61936 62140 62000
rect 62204 61936 62220 62000
rect 62284 61936 62322 62000
rect 61702 52240 62322 61936
rect 61702 52176 61740 52240
rect 61804 52176 61820 52240
rect 61884 52176 61900 52240
rect 61964 52176 61980 52240
rect 62044 52176 62060 52240
rect 62124 52176 62140 52240
rect 62204 52176 62220 52240
rect 62284 52176 62322 52240
rect 61702 52160 62322 52176
rect 61702 52096 61740 52160
rect 61804 52096 61820 52160
rect 61884 52096 61900 52160
rect 61964 52096 61980 52160
rect 62044 52096 62060 52160
rect 62124 52096 62140 52160
rect 62204 52096 62220 52160
rect 62284 52096 62322 52160
rect 61702 52080 62322 52096
rect 61702 52016 61740 52080
rect 61804 52016 61820 52080
rect 61884 52016 61900 52080
rect 61964 52016 61980 52080
rect 62044 52016 62060 52080
rect 62124 52016 62140 52080
rect 62204 52016 62220 52080
rect 62284 52016 62322 52080
rect 61702 52000 62322 52016
rect 61702 51936 61740 52000
rect 61804 51936 61820 52000
rect 61884 51936 61900 52000
rect 61964 51936 61980 52000
rect 62044 51936 62060 52000
rect 62124 51936 62140 52000
rect 62204 51936 62220 52000
rect 62284 51936 62322 52000
rect 61702 42240 62322 51936
rect 61702 42176 61740 42240
rect 61804 42176 61820 42240
rect 61884 42176 61900 42240
rect 61964 42176 61980 42240
rect 62044 42176 62060 42240
rect 62124 42176 62140 42240
rect 62204 42176 62220 42240
rect 62284 42176 62322 42240
rect 61702 42160 62322 42176
rect 61702 42096 61740 42160
rect 61804 42096 61820 42160
rect 61884 42096 61900 42160
rect 61964 42096 61980 42160
rect 62044 42096 62060 42160
rect 62124 42096 62140 42160
rect 62204 42096 62220 42160
rect 62284 42096 62322 42160
rect 61702 42080 62322 42096
rect 61702 42016 61740 42080
rect 61804 42016 61820 42080
rect 61884 42016 61900 42080
rect 61964 42016 61980 42080
rect 62044 42016 62060 42080
rect 62124 42016 62140 42080
rect 62204 42016 62220 42080
rect 62284 42016 62322 42080
rect 61702 42000 62322 42016
rect 61702 41936 61740 42000
rect 61804 41936 61820 42000
rect 61884 41936 61900 42000
rect 61964 41936 61980 42000
rect 62044 41936 62060 42000
rect 62124 41936 62140 42000
rect 62204 41936 62220 42000
rect 62284 41936 62322 42000
rect 61702 32240 62322 41936
rect 61702 32176 61740 32240
rect 61804 32176 61820 32240
rect 61884 32176 61900 32240
rect 61964 32176 61980 32240
rect 62044 32176 62060 32240
rect 62124 32176 62140 32240
rect 62204 32176 62220 32240
rect 62284 32176 62322 32240
rect 61702 32160 62322 32176
rect 61702 32096 61740 32160
rect 61804 32096 61820 32160
rect 61884 32096 61900 32160
rect 61964 32096 61980 32160
rect 62044 32096 62060 32160
rect 62124 32096 62140 32160
rect 62204 32096 62220 32160
rect 62284 32096 62322 32160
rect 61702 32080 62322 32096
rect 61702 32016 61740 32080
rect 61804 32016 61820 32080
rect 61884 32016 61900 32080
rect 61964 32016 61980 32080
rect 62044 32016 62060 32080
rect 62124 32016 62140 32080
rect 62204 32016 62220 32080
rect 62284 32016 62322 32080
rect 61702 32000 62322 32016
rect 61702 31936 61740 32000
rect 61804 31936 61820 32000
rect 61884 31936 61900 32000
rect 61964 31936 61980 32000
rect 62044 31936 62060 32000
rect 62124 31936 62140 32000
rect 62204 31936 62220 32000
rect 62284 31936 62322 32000
rect 61702 22240 62322 31936
rect 61702 22176 61740 22240
rect 61804 22176 61820 22240
rect 61884 22176 61900 22240
rect 61964 22176 61980 22240
rect 62044 22176 62060 22240
rect 62124 22176 62140 22240
rect 62204 22176 62220 22240
rect 62284 22176 62322 22240
rect 61702 22160 62322 22176
rect 61702 22096 61740 22160
rect 61804 22096 61820 22160
rect 61884 22096 61900 22160
rect 61964 22096 61980 22160
rect 62044 22096 62060 22160
rect 62124 22096 62140 22160
rect 62204 22096 62220 22160
rect 62284 22096 62322 22160
rect 61702 22080 62322 22096
rect 61702 22016 61740 22080
rect 61804 22016 61820 22080
rect 61884 22016 61900 22080
rect 61964 22016 61980 22080
rect 62044 22016 62060 22080
rect 62124 22016 62140 22080
rect 62204 22016 62220 22080
rect 62284 22016 62322 22080
rect 61702 22000 62322 22016
rect 61702 21936 61740 22000
rect 61804 21936 61820 22000
rect 61884 21936 61900 22000
rect 61964 21936 61980 22000
rect 62044 21936 62060 22000
rect 62124 21936 62140 22000
rect 62204 21936 62220 22000
rect 62284 21936 62322 22000
rect 61702 12240 62322 21936
rect 63171 15876 63237 15877
rect 63171 15812 63172 15876
rect 63236 15812 63237 15876
rect 63171 15811 63237 15812
rect 61702 12176 61740 12240
rect 61804 12176 61820 12240
rect 61884 12176 61900 12240
rect 61964 12176 61980 12240
rect 62044 12176 62060 12240
rect 62124 12176 62140 12240
rect 62204 12176 62220 12240
rect 62284 12176 62322 12240
rect 61702 12160 62322 12176
rect 61702 12096 61740 12160
rect 61804 12096 61820 12160
rect 61884 12096 61900 12160
rect 61964 12096 61980 12160
rect 62044 12096 62060 12160
rect 62124 12096 62140 12160
rect 62204 12096 62220 12160
rect 62284 12096 62322 12160
rect 61702 12080 62322 12096
rect 61702 12016 61740 12080
rect 61804 12016 61820 12080
rect 61884 12016 61900 12080
rect 61964 12016 61980 12080
rect 62044 12016 62060 12080
rect 62124 12016 62140 12080
rect 62204 12016 62220 12080
rect 62284 12016 62322 12080
rect 61702 12000 62322 12016
rect 61702 11936 61740 12000
rect 61804 11936 61820 12000
rect 61884 11936 61900 12000
rect 61964 11936 61980 12000
rect 62044 11936 62060 12000
rect 62124 11936 62140 12000
rect 62204 11936 62220 12000
rect 62284 11936 62322 12000
rect 61702 2240 62322 11936
rect 62987 10572 63053 10573
rect 62987 10508 62988 10572
rect 63052 10508 63053 10572
rect 62987 10507 63053 10508
rect 62990 7173 63050 10507
rect 63174 9893 63234 15811
rect 63355 11524 63421 11525
rect 63355 11460 63356 11524
rect 63420 11460 63421 11524
rect 63355 11459 63421 11460
rect 63358 10029 63418 11459
rect 63355 10028 63421 10029
rect 63355 9964 63356 10028
rect 63420 9964 63421 10028
rect 63355 9963 63421 9964
rect 63171 9892 63237 9893
rect 63171 9828 63172 9892
rect 63236 9828 63237 9892
rect 63171 9827 63237 9828
rect 62987 7172 63053 7173
rect 62987 7108 62988 7172
rect 63052 7108 63053 7172
rect 62987 7107 63053 7108
rect 63358 5541 63418 9963
rect 63542 7581 63602 65179
rect 64702 64592 65322 74288
rect 64702 64528 64740 64592
rect 64804 64528 64820 64592
rect 64884 64528 64900 64592
rect 64964 64528 64980 64592
rect 65044 64528 65060 64592
rect 65124 64528 65140 64592
rect 65204 64528 65220 64592
rect 65284 64528 65322 64592
rect 64702 64512 65322 64528
rect 64702 64448 64740 64512
rect 64804 64448 64820 64512
rect 64884 64448 64900 64512
rect 64964 64448 64980 64512
rect 65044 64448 65060 64512
rect 65124 64448 65140 64512
rect 65204 64448 65220 64512
rect 65284 64448 65322 64512
rect 64702 64432 65322 64448
rect 64702 64368 64740 64432
rect 64804 64368 64820 64432
rect 64884 64368 64900 64432
rect 64964 64368 64980 64432
rect 65044 64368 65060 64432
rect 65124 64368 65140 64432
rect 65204 64368 65220 64432
rect 65284 64368 65322 64432
rect 64702 64352 65322 64368
rect 64702 64288 64740 64352
rect 64804 64288 64820 64352
rect 64884 64288 64900 64352
rect 64964 64288 64980 64352
rect 65044 64288 65060 64352
rect 65124 64288 65140 64352
rect 65204 64288 65220 64352
rect 65284 64288 65322 64352
rect 63723 63204 63789 63205
rect 63723 63140 63724 63204
rect 63788 63140 63789 63204
rect 63723 63139 63789 63140
rect 63539 7580 63605 7581
rect 63539 7516 63540 7580
rect 63604 7516 63605 7580
rect 63539 7515 63605 7516
rect 63726 5949 63786 63139
rect 63907 61028 63973 61029
rect 63907 60964 63908 61028
rect 63972 60964 63973 61028
rect 63907 60963 63973 60964
rect 63910 6765 63970 60963
rect 64091 58716 64157 58717
rect 64091 58652 64092 58716
rect 64156 58652 64157 58716
rect 64091 58651 64157 58652
rect 63907 6764 63973 6765
rect 63907 6700 63908 6764
rect 63972 6700 63973 6764
rect 63907 6699 63973 6700
rect 63723 5948 63789 5949
rect 63723 5884 63724 5948
rect 63788 5884 63789 5948
rect 63723 5883 63789 5884
rect 63355 5540 63421 5541
rect 63355 5476 63356 5540
rect 63420 5476 63421 5540
rect 63355 5475 63421 5476
rect 64094 3365 64154 58651
rect 64275 56676 64341 56677
rect 64275 56612 64276 56676
rect 64340 56612 64341 56676
rect 64275 56611 64341 56612
rect 64278 6629 64338 56611
rect 64702 54592 65322 64288
rect 64702 54528 64740 54592
rect 64804 54528 64820 54592
rect 64884 54528 64900 54592
rect 64964 54528 64980 54592
rect 65044 54528 65060 54592
rect 65124 54528 65140 54592
rect 65204 54528 65220 54592
rect 65284 54528 65322 54592
rect 64702 54512 65322 54528
rect 64702 54448 64740 54512
rect 64804 54448 64820 54512
rect 64884 54448 64900 54512
rect 64964 54448 64980 54512
rect 65044 54448 65060 54512
rect 65124 54448 65140 54512
rect 65204 54448 65220 54512
rect 65284 54448 65322 54512
rect 64702 54432 65322 54448
rect 64702 54368 64740 54432
rect 64804 54368 64820 54432
rect 64884 54368 64900 54432
rect 64964 54368 64980 54432
rect 65044 54368 65060 54432
rect 65124 54368 65140 54432
rect 65204 54368 65220 54432
rect 65284 54368 65322 54432
rect 64702 54352 65322 54368
rect 64702 54288 64740 54352
rect 64804 54288 64820 54352
rect 64884 54288 64900 54352
rect 64964 54288 64980 54352
rect 65044 54288 65060 54352
rect 65124 54288 65140 54352
rect 65204 54288 65220 54352
rect 65284 54288 65322 54352
rect 64702 44592 65322 54288
rect 67702 82240 68322 87000
rect 67702 82176 67740 82240
rect 67804 82176 67820 82240
rect 67884 82176 67900 82240
rect 67964 82176 67980 82240
rect 68044 82176 68060 82240
rect 68124 82176 68140 82240
rect 68204 82176 68220 82240
rect 68284 82176 68322 82240
rect 67702 82160 68322 82176
rect 67702 82096 67740 82160
rect 67804 82096 67820 82160
rect 67884 82096 67900 82160
rect 67964 82096 67980 82160
rect 68044 82096 68060 82160
rect 68124 82096 68140 82160
rect 68204 82096 68220 82160
rect 68284 82096 68322 82160
rect 67702 82080 68322 82096
rect 67702 82016 67740 82080
rect 67804 82016 67820 82080
rect 67884 82016 67900 82080
rect 67964 82016 67980 82080
rect 68044 82016 68060 82080
rect 68124 82016 68140 82080
rect 68204 82016 68220 82080
rect 68284 82016 68322 82080
rect 67702 82000 68322 82016
rect 67702 81936 67740 82000
rect 67804 81936 67820 82000
rect 67884 81936 67900 82000
rect 67964 81936 67980 82000
rect 68044 81936 68060 82000
rect 68124 81936 68140 82000
rect 68204 81936 68220 82000
rect 68284 81936 68322 82000
rect 67702 72240 68322 81936
rect 67702 72176 67740 72240
rect 67804 72176 67820 72240
rect 67884 72176 67900 72240
rect 67964 72176 67980 72240
rect 68044 72176 68060 72240
rect 68124 72176 68140 72240
rect 68204 72176 68220 72240
rect 68284 72176 68322 72240
rect 67702 72160 68322 72176
rect 67702 72096 67740 72160
rect 67804 72096 67820 72160
rect 67884 72096 67900 72160
rect 67964 72096 67980 72160
rect 68044 72096 68060 72160
rect 68124 72096 68140 72160
rect 68204 72096 68220 72160
rect 68284 72096 68322 72160
rect 67702 72080 68322 72096
rect 67702 72016 67740 72080
rect 67804 72016 67820 72080
rect 67884 72016 67900 72080
rect 67964 72016 67980 72080
rect 68044 72016 68060 72080
rect 68124 72016 68140 72080
rect 68204 72016 68220 72080
rect 68284 72016 68322 72080
rect 67702 72000 68322 72016
rect 67702 71936 67740 72000
rect 67804 71936 67820 72000
rect 67884 71936 67900 72000
rect 67964 71936 67980 72000
rect 68044 71936 68060 72000
rect 68124 71936 68140 72000
rect 68204 71936 68220 72000
rect 68284 71936 68322 72000
rect 67702 62240 68322 71936
rect 67702 62176 67740 62240
rect 67804 62176 67820 62240
rect 67884 62176 67900 62240
rect 67964 62176 67980 62240
rect 68044 62176 68060 62240
rect 68124 62176 68140 62240
rect 68204 62176 68220 62240
rect 68284 62176 68322 62240
rect 67702 62160 68322 62176
rect 67702 62096 67740 62160
rect 67804 62096 67820 62160
rect 67884 62096 67900 62160
rect 67964 62096 67980 62160
rect 68044 62096 68060 62160
rect 68124 62096 68140 62160
rect 68204 62096 68220 62160
rect 68284 62096 68322 62160
rect 67702 62080 68322 62096
rect 67702 62016 67740 62080
rect 67804 62016 67820 62080
rect 67884 62016 67900 62080
rect 67964 62016 67980 62080
rect 68044 62016 68060 62080
rect 68124 62016 68140 62080
rect 68204 62016 68220 62080
rect 68284 62016 68322 62080
rect 67702 62000 68322 62016
rect 67702 61936 67740 62000
rect 67804 61936 67820 62000
rect 67884 61936 67900 62000
rect 67964 61936 67980 62000
rect 68044 61936 68060 62000
rect 68124 61936 68140 62000
rect 68204 61936 68220 62000
rect 68284 61936 68322 62000
rect 67702 52240 68322 61936
rect 70702 84592 71322 87000
rect 70702 84528 70740 84592
rect 70804 84528 70820 84592
rect 70884 84528 70900 84592
rect 70964 84528 70980 84592
rect 71044 84528 71060 84592
rect 71124 84528 71140 84592
rect 71204 84528 71220 84592
rect 71284 84528 71322 84592
rect 70702 84512 71322 84528
rect 70702 84448 70740 84512
rect 70804 84448 70820 84512
rect 70884 84448 70900 84512
rect 70964 84448 70980 84512
rect 71044 84448 71060 84512
rect 71124 84448 71140 84512
rect 71204 84448 71220 84512
rect 71284 84448 71322 84512
rect 70702 84432 71322 84448
rect 70702 84368 70740 84432
rect 70804 84368 70820 84432
rect 70884 84368 70900 84432
rect 70964 84368 70980 84432
rect 71044 84368 71060 84432
rect 71124 84368 71140 84432
rect 71204 84368 71220 84432
rect 71284 84368 71322 84432
rect 70702 84352 71322 84368
rect 70702 84288 70740 84352
rect 70804 84288 70820 84352
rect 70884 84288 70900 84352
rect 70964 84288 70980 84352
rect 71044 84288 71060 84352
rect 71124 84288 71140 84352
rect 71204 84288 71220 84352
rect 71284 84288 71322 84352
rect 70702 74592 71322 84288
rect 70702 74528 70740 74592
rect 70804 74528 70820 74592
rect 70884 74528 70900 74592
rect 70964 74528 70980 74592
rect 71044 74528 71060 74592
rect 71124 74528 71140 74592
rect 71204 74528 71220 74592
rect 71284 74528 71322 74592
rect 70702 74512 71322 74528
rect 70702 74448 70740 74512
rect 70804 74448 70820 74512
rect 70884 74448 70900 74512
rect 70964 74448 70980 74512
rect 71044 74448 71060 74512
rect 71124 74448 71140 74512
rect 71204 74448 71220 74512
rect 71284 74448 71322 74512
rect 70702 74432 71322 74448
rect 70702 74368 70740 74432
rect 70804 74368 70820 74432
rect 70884 74368 70900 74432
rect 70964 74368 70980 74432
rect 71044 74368 71060 74432
rect 71124 74368 71140 74432
rect 71204 74368 71220 74432
rect 71284 74368 71322 74432
rect 70702 74352 71322 74368
rect 70702 74288 70740 74352
rect 70804 74288 70820 74352
rect 70884 74288 70900 74352
rect 70964 74288 70980 74352
rect 71044 74288 71060 74352
rect 71124 74288 71140 74352
rect 71204 74288 71220 74352
rect 71284 74288 71322 74352
rect 70702 64592 71322 74288
rect 70702 64528 70740 64592
rect 70804 64528 70820 64592
rect 70884 64528 70900 64592
rect 70964 64528 70980 64592
rect 71044 64528 71060 64592
rect 71124 64528 71140 64592
rect 71204 64528 71220 64592
rect 71284 64528 71322 64592
rect 70702 64512 71322 64528
rect 70702 64448 70740 64512
rect 70804 64448 70820 64512
rect 70884 64448 70900 64512
rect 70964 64448 70980 64512
rect 71044 64448 71060 64512
rect 71124 64448 71140 64512
rect 71204 64448 71220 64512
rect 71284 64448 71322 64512
rect 70702 64432 71322 64448
rect 70702 64368 70740 64432
rect 70804 64368 70820 64432
rect 70884 64368 70900 64432
rect 70964 64368 70980 64432
rect 71044 64368 71060 64432
rect 71124 64368 71140 64432
rect 71204 64368 71220 64432
rect 71284 64368 71322 64432
rect 70702 64352 71322 64368
rect 70702 64288 70740 64352
rect 70804 64288 70820 64352
rect 70884 64288 70900 64352
rect 70964 64288 70980 64352
rect 71044 64288 71060 64352
rect 71124 64288 71140 64352
rect 71204 64288 71220 64352
rect 71284 64288 71322 64352
rect 69059 54772 69125 54773
rect 69059 54708 69060 54772
rect 69124 54708 69125 54772
rect 69059 54707 69125 54708
rect 67702 52176 67740 52240
rect 67804 52176 67820 52240
rect 67884 52176 67900 52240
rect 67964 52176 67980 52240
rect 68044 52176 68060 52240
rect 68124 52176 68140 52240
rect 68204 52176 68220 52240
rect 68284 52176 68322 52240
rect 67702 52160 68322 52176
rect 67702 52096 67740 52160
rect 67804 52096 67820 52160
rect 67884 52096 67900 52160
rect 67964 52096 67980 52160
rect 68044 52096 68060 52160
rect 68124 52096 68140 52160
rect 68204 52096 68220 52160
rect 68284 52096 68322 52160
rect 67702 52080 68322 52096
rect 67702 52016 67740 52080
rect 67804 52016 67820 52080
rect 67884 52016 67900 52080
rect 67964 52016 67980 52080
rect 68044 52016 68060 52080
rect 68124 52016 68140 52080
rect 68204 52016 68220 52080
rect 68284 52016 68322 52080
rect 67702 52000 68322 52016
rect 67702 51936 67740 52000
rect 67804 51936 67820 52000
rect 67884 51936 67900 52000
rect 67964 51936 67980 52000
rect 68044 51936 68060 52000
rect 68124 51936 68140 52000
rect 68204 51936 68220 52000
rect 68284 51936 68322 52000
rect 65747 47020 65813 47021
rect 65747 46956 65748 47020
rect 65812 46956 65813 47020
rect 65747 46955 65813 46956
rect 66115 47020 66181 47021
rect 66115 46956 66116 47020
rect 66180 46956 66181 47020
rect 66115 46955 66181 46956
rect 64702 44528 64740 44592
rect 64804 44528 64820 44592
rect 64884 44528 64900 44592
rect 64964 44528 64980 44592
rect 65044 44528 65060 44592
rect 65124 44528 65140 44592
rect 65204 44528 65220 44592
rect 65284 44528 65322 44592
rect 64702 44512 65322 44528
rect 64702 44448 64740 44512
rect 64804 44448 64820 44512
rect 64884 44448 64900 44512
rect 64964 44448 64980 44512
rect 65044 44448 65060 44512
rect 65124 44448 65140 44512
rect 65204 44448 65220 44512
rect 65284 44448 65322 44512
rect 64702 44432 65322 44448
rect 64702 44368 64740 44432
rect 64804 44368 64820 44432
rect 64884 44368 64900 44432
rect 64964 44368 64980 44432
rect 65044 44368 65060 44432
rect 65124 44368 65140 44432
rect 65204 44368 65220 44432
rect 65284 44368 65322 44432
rect 64702 44352 65322 44368
rect 64702 44288 64740 44352
rect 64804 44288 64820 44352
rect 64884 44288 64900 44352
rect 64964 44288 64980 44352
rect 65044 44288 65060 44352
rect 65124 44288 65140 44352
rect 65204 44288 65220 44352
rect 65284 44288 65322 44352
rect 64702 34592 65322 44288
rect 65563 41308 65629 41309
rect 65563 41244 65564 41308
rect 65628 41244 65629 41308
rect 65563 41243 65629 41244
rect 65566 38589 65626 41243
rect 65563 38588 65629 38589
rect 65563 38524 65564 38588
rect 65628 38524 65629 38588
rect 65563 38523 65629 38524
rect 65563 34780 65629 34781
rect 65563 34716 65564 34780
rect 65628 34716 65629 34780
rect 65563 34715 65629 34716
rect 64702 34528 64740 34592
rect 64804 34528 64820 34592
rect 64884 34528 64900 34592
rect 64964 34528 64980 34592
rect 65044 34528 65060 34592
rect 65124 34528 65140 34592
rect 65204 34528 65220 34592
rect 65284 34528 65322 34592
rect 64702 34512 65322 34528
rect 64702 34448 64740 34512
rect 64804 34448 64820 34512
rect 64884 34448 64900 34512
rect 64964 34448 64980 34512
rect 65044 34448 65060 34512
rect 65124 34448 65140 34512
rect 65204 34448 65220 34512
rect 65284 34448 65322 34512
rect 64702 34432 65322 34448
rect 64702 34368 64740 34432
rect 64804 34368 64820 34432
rect 64884 34368 64900 34432
rect 64964 34368 64980 34432
rect 65044 34368 65060 34432
rect 65124 34368 65140 34432
rect 65204 34368 65220 34432
rect 65284 34368 65322 34432
rect 64702 34352 65322 34368
rect 64702 34288 64740 34352
rect 64804 34288 64820 34352
rect 64884 34288 64900 34352
rect 64964 34288 64980 34352
rect 65044 34288 65060 34352
rect 65124 34288 65140 34352
rect 65204 34288 65220 34352
rect 65284 34288 65322 34352
rect 64702 24592 65322 34288
rect 64702 24528 64740 24592
rect 64804 24528 64820 24592
rect 64884 24528 64900 24592
rect 64964 24528 64980 24592
rect 65044 24528 65060 24592
rect 65124 24528 65140 24592
rect 65204 24528 65220 24592
rect 65284 24528 65322 24592
rect 64702 24512 65322 24528
rect 64702 24448 64740 24512
rect 64804 24448 64820 24512
rect 64884 24448 64900 24512
rect 64964 24448 64980 24512
rect 65044 24448 65060 24512
rect 65124 24448 65140 24512
rect 65204 24448 65220 24512
rect 65284 24448 65322 24512
rect 64702 24432 65322 24448
rect 64702 24368 64740 24432
rect 64804 24368 64820 24432
rect 64884 24368 64900 24432
rect 64964 24368 64980 24432
rect 65044 24368 65060 24432
rect 65124 24368 65140 24432
rect 65204 24368 65220 24432
rect 65284 24368 65322 24432
rect 64702 24352 65322 24368
rect 64702 24288 64740 24352
rect 64804 24288 64820 24352
rect 64884 24288 64900 24352
rect 64964 24288 64980 24352
rect 65044 24288 65060 24352
rect 65124 24288 65140 24352
rect 65204 24288 65220 24352
rect 65284 24288 65322 24352
rect 64459 18188 64525 18189
rect 64459 18124 64460 18188
rect 64524 18124 64525 18188
rect 64459 18123 64525 18124
rect 64462 11797 64522 18123
rect 64702 14592 65322 24288
rect 64702 14528 64740 14592
rect 64804 14528 64820 14592
rect 64884 14528 64900 14592
rect 64964 14528 64980 14592
rect 65044 14528 65060 14592
rect 65124 14528 65140 14592
rect 65204 14528 65220 14592
rect 65284 14528 65322 14592
rect 64702 14512 65322 14528
rect 64702 14448 64740 14512
rect 64804 14448 64820 14512
rect 64884 14448 64900 14512
rect 64964 14448 64980 14512
rect 65044 14448 65060 14512
rect 65124 14448 65140 14512
rect 65204 14448 65220 14512
rect 65284 14448 65322 14512
rect 64702 14432 65322 14448
rect 64702 14368 64740 14432
rect 64804 14368 64820 14432
rect 64884 14368 64900 14432
rect 64964 14368 64980 14432
rect 65044 14368 65060 14432
rect 65124 14368 65140 14432
rect 65204 14368 65220 14432
rect 65284 14368 65322 14432
rect 64702 14352 65322 14368
rect 64702 14288 64740 14352
rect 64804 14288 64820 14352
rect 64884 14288 64900 14352
rect 64964 14288 64980 14352
rect 65044 14288 65060 14352
rect 65124 14288 65140 14352
rect 65204 14288 65220 14352
rect 65284 14288 65322 14352
rect 64459 11796 64525 11797
rect 64459 11732 64460 11796
rect 64524 11732 64525 11796
rect 64459 11731 64525 11732
rect 64275 6628 64341 6629
rect 64275 6564 64276 6628
rect 64340 6564 64341 6628
rect 64275 6563 64341 6564
rect 64702 4592 65322 14288
rect 64702 4528 64740 4592
rect 64804 4528 64820 4592
rect 64884 4528 64900 4592
rect 64964 4528 64980 4592
rect 65044 4528 65060 4592
rect 65124 4528 65140 4592
rect 65204 4528 65220 4592
rect 65284 4528 65322 4592
rect 64702 4512 65322 4528
rect 64702 4448 64740 4512
rect 64804 4448 64820 4512
rect 64884 4448 64900 4512
rect 64964 4448 64980 4512
rect 65044 4448 65060 4512
rect 65124 4448 65140 4512
rect 65204 4448 65220 4512
rect 65284 4448 65322 4512
rect 64702 4432 65322 4448
rect 64702 4368 64740 4432
rect 64804 4368 64820 4432
rect 64884 4368 64900 4432
rect 64964 4368 64980 4432
rect 65044 4368 65060 4432
rect 65124 4368 65140 4432
rect 65204 4368 65220 4432
rect 65284 4368 65322 4432
rect 64702 4352 65322 4368
rect 64702 4288 64740 4352
rect 64804 4288 64820 4352
rect 64884 4288 64900 4352
rect 64964 4288 64980 4352
rect 65044 4288 65060 4352
rect 65124 4288 65140 4352
rect 65204 4288 65220 4352
rect 65284 4288 65322 4352
rect 64091 3364 64157 3365
rect 64091 3300 64092 3364
rect 64156 3300 64157 3364
rect 64091 3299 64157 3300
rect 61702 2176 61740 2240
rect 61804 2176 61820 2240
rect 61884 2176 61900 2240
rect 61964 2176 61980 2240
rect 62044 2176 62060 2240
rect 62124 2176 62140 2240
rect 62204 2176 62220 2240
rect 62284 2176 62322 2240
rect 61702 2160 62322 2176
rect 61702 2096 61740 2160
rect 61804 2096 61820 2160
rect 61884 2096 61900 2160
rect 61964 2096 61980 2160
rect 62044 2096 62060 2160
rect 62124 2096 62140 2160
rect 62204 2096 62220 2160
rect 62284 2096 62322 2160
rect 61702 2080 62322 2096
rect 61702 2016 61740 2080
rect 61804 2016 61820 2080
rect 61884 2016 61900 2080
rect 61964 2016 61980 2080
rect 62044 2016 62060 2080
rect 62124 2016 62140 2080
rect 62204 2016 62220 2080
rect 62284 2016 62322 2080
rect 61702 2000 62322 2016
rect 61702 1936 61740 2000
rect 61804 1936 61820 2000
rect 61884 1936 61900 2000
rect 61964 1936 61980 2000
rect 62044 1936 62060 2000
rect 62124 1936 62140 2000
rect 62204 1936 62220 2000
rect 62284 1936 62322 2000
rect 61702 0 62322 1936
rect 64702 0 65322 4288
rect 65566 1325 65626 34715
rect 65750 7853 65810 46955
rect 65931 12748 65997 12749
rect 65931 12684 65932 12748
rect 65996 12684 65997 12748
rect 65931 12683 65997 12684
rect 65934 11797 65994 12683
rect 65931 11796 65997 11797
rect 65931 11732 65932 11796
rect 65996 11732 65997 11796
rect 65931 11731 65997 11732
rect 65747 7852 65813 7853
rect 65747 7788 65748 7852
rect 65812 7788 65813 7852
rect 65747 7787 65813 7788
rect 66118 7445 66178 46955
rect 67702 42240 68322 51936
rect 67702 42176 67740 42240
rect 67804 42176 67820 42240
rect 67884 42176 67900 42240
rect 67964 42176 67980 42240
rect 68044 42176 68060 42240
rect 68124 42176 68140 42240
rect 68204 42176 68220 42240
rect 68284 42176 68322 42240
rect 67702 42160 68322 42176
rect 67702 42096 67740 42160
rect 67804 42096 67820 42160
rect 67884 42096 67900 42160
rect 67964 42096 67980 42160
rect 68044 42096 68060 42160
rect 68124 42096 68140 42160
rect 68204 42096 68220 42160
rect 68284 42096 68322 42160
rect 67702 42080 68322 42096
rect 67702 42016 67740 42080
rect 67804 42016 67820 42080
rect 67884 42016 67900 42080
rect 67964 42016 67980 42080
rect 68044 42016 68060 42080
rect 68124 42016 68140 42080
rect 68204 42016 68220 42080
rect 68284 42016 68322 42080
rect 67702 42000 68322 42016
rect 67702 41936 67740 42000
rect 67804 41936 67820 42000
rect 67884 41936 67900 42000
rect 67964 41936 67980 42000
rect 68044 41936 68060 42000
rect 68124 41936 68140 42000
rect 68204 41936 68220 42000
rect 68284 41936 68322 42000
rect 67702 32240 68322 41936
rect 67702 32176 67740 32240
rect 67804 32176 67820 32240
rect 67884 32176 67900 32240
rect 67964 32176 67980 32240
rect 68044 32176 68060 32240
rect 68124 32176 68140 32240
rect 68204 32176 68220 32240
rect 68284 32176 68322 32240
rect 67702 32160 68322 32176
rect 67702 32096 67740 32160
rect 67804 32096 67820 32160
rect 67884 32096 67900 32160
rect 67964 32096 67980 32160
rect 68044 32096 68060 32160
rect 68124 32096 68140 32160
rect 68204 32096 68220 32160
rect 68284 32096 68322 32160
rect 67702 32080 68322 32096
rect 67702 32016 67740 32080
rect 67804 32016 67820 32080
rect 67884 32016 67900 32080
rect 67964 32016 67980 32080
rect 68044 32016 68060 32080
rect 68124 32016 68140 32080
rect 68204 32016 68220 32080
rect 68284 32016 68322 32080
rect 67702 32000 68322 32016
rect 67702 31936 67740 32000
rect 67804 31936 67820 32000
rect 67884 31936 67900 32000
rect 67964 31936 67980 32000
rect 68044 31936 68060 32000
rect 68124 31936 68140 32000
rect 68204 31936 68220 32000
rect 68284 31936 68322 32000
rect 67035 23628 67101 23629
rect 67035 23564 67036 23628
rect 67100 23564 67101 23628
rect 67035 23563 67101 23564
rect 66483 22676 66549 22677
rect 66483 22612 66484 22676
rect 66548 22612 66549 22676
rect 66483 22611 66549 22612
rect 66299 22404 66365 22405
rect 66299 22340 66300 22404
rect 66364 22340 66365 22404
rect 66299 22339 66365 22340
rect 66115 7444 66181 7445
rect 66115 7380 66116 7444
rect 66180 7380 66181 7444
rect 66115 7379 66181 7380
rect 66302 7037 66362 22339
rect 66299 7036 66365 7037
rect 66299 6972 66300 7036
rect 66364 6972 66365 7036
rect 66299 6971 66365 6972
rect 66486 3909 66546 22611
rect 67038 7309 67098 23563
rect 67219 23492 67285 23493
rect 67219 23428 67220 23492
rect 67284 23428 67285 23492
rect 67219 23427 67285 23428
rect 67035 7308 67101 7309
rect 67035 7244 67036 7308
rect 67100 7244 67101 7308
rect 67035 7243 67101 7244
rect 66483 3908 66549 3909
rect 66483 3844 66484 3908
rect 66548 3844 66549 3908
rect 66483 3843 66549 3844
rect 67222 3093 67282 23427
rect 67702 22240 68322 31936
rect 67702 22176 67740 22240
rect 67804 22176 67820 22240
rect 67884 22176 67900 22240
rect 67964 22176 67980 22240
rect 68044 22176 68060 22240
rect 68124 22176 68140 22240
rect 68204 22176 68220 22240
rect 68284 22176 68322 22240
rect 67702 22160 68322 22176
rect 67702 22096 67740 22160
rect 67804 22096 67820 22160
rect 67884 22096 67900 22160
rect 67964 22096 67980 22160
rect 68044 22096 68060 22160
rect 68124 22096 68140 22160
rect 68204 22096 68220 22160
rect 68284 22096 68322 22160
rect 67702 22080 68322 22096
rect 67702 22016 67740 22080
rect 67804 22016 67820 22080
rect 67884 22016 67900 22080
rect 67964 22016 67980 22080
rect 68044 22016 68060 22080
rect 68124 22016 68140 22080
rect 68204 22016 68220 22080
rect 68284 22016 68322 22080
rect 67702 22000 68322 22016
rect 67702 21936 67740 22000
rect 67804 21936 67820 22000
rect 67884 21936 67900 22000
rect 67964 21936 67980 22000
rect 68044 21936 68060 22000
rect 68124 21936 68140 22000
rect 68204 21936 68220 22000
rect 68284 21936 68322 22000
rect 67702 12240 68322 21936
rect 67702 12176 67740 12240
rect 67804 12176 67820 12240
rect 67884 12176 67900 12240
rect 67964 12176 67980 12240
rect 68044 12176 68060 12240
rect 68124 12176 68140 12240
rect 68204 12176 68220 12240
rect 68284 12176 68322 12240
rect 67702 12160 68322 12176
rect 67702 12096 67740 12160
rect 67804 12096 67820 12160
rect 67884 12096 67900 12160
rect 67964 12096 67980 12160
rect 68044 12096 68060 12160
rect 68124 12096 68140 12160
rect 68204 12096 68220 12160
rect 68284 12096 68322 12160
rect 67702 12080 68322 12096
rect 67702 12016 67740 12080
rect 67804 12016 67820 12080
rect 67884 12016 67900 12080
rect 67964 12016 67980 12080
rect 68044 12016 68060 12080
rect 68124 12016 68140 12080
rect 68204 12016 68220 12080
rect 68284 12016 68322 12080
rect 67702 12000 68322 12016
rect 67702 11936 67740 12000
rect 67804 11936 67820 12000
rect 67884 11936 67900 12000
rect 67964 11936 67980 12000
rect 68044 11936 68060 12000
rect 68124 11936 68140 12000
rect 68204 11936 68220 12000
rect 68284 11936 68322 12000
rect 67219 3092 67285 3093
rect 67219 3028 67220 3092
rect 67284 3028 67285 3092
rect 67219 3027 67285 3028
rect 67702 2240 68322 11936
rect 69062 3773 69122 54707
rect 70702 54592 71322 64288
rect 70702 54528 70740 54592
rect 70804 54528 70820 54592
rect 70884 54528 70900 54592
rect 70964 54528 70980 54592
rect 71044 54528 71060 54592
rect 71124 54528 71140 54592
rect 71204 54528 71220 54592
rect 71284 54528 71322 54592
rect 70702 54512 71322 54528
rect 70702 54448 70740 54512
rect 70804 54448 70820 54512
rect 70884 54448 70900 54512
rect 70964 54448 70980 54512
rect 71044 54448 71060 54512
rect 71124 54448 71140 54512
rect 71204 54448 71220 54512
rect 71284 54448 71322 54512
rect 70702 54432 71322 54448
rect 70702 54368 70740 54432
rect 70804 54368 70820 54432
rect 70884 54368 70900 54432
rect 70964 54368 70980 54432
rect 71044 54368 71060 54432
rect 71124 54368 71140 54432
rect 71204 54368 71220 54432
rect 71284 54368 71322 54432
rect 70702 54352 71322 54368
rect 70702 54288 70740 54352
rect 70804 54288 70820 54352
rect 70884 54288 70900 54352
rect 70964 54288 70980 54352
rect 71044 54288 71060 54352
rect 71124 54288 71140 54352
rect 71204 54288 71220 54352
rect 71284 54288 71322 54352
rect 70702 44592 71322 54288
rect 70702 44528 70740 44592
rect 70804 44528 70820 44592
rect 70884 44528 70900 44592
rect 70964 44528 70980 44592
rect 71044 44528 71060 44592
rect 71124 44528 71140 44592
rect 71204 44528 71220 44592
rect 71284 44528 71322 44592
rect 70702 44512 71322 44528
rect 70702 44448 70740 44512
rect 70804 44448 70820 44512
rect 70884 44448 70900 44512
rect 70964 44448 70980 44512
rect 71044 44448 71060 44512
rect 71124 44448 71140 44512
rect 71204 44448 71220 44512
rect 71284 44448 71322 44512
rect 70702 44432 71322 44448
rect 70702 44368 70740 44432
rect 70804 44368 70820 44432
rect 70884 44368 70900 44432
rect 70964 44368 70980 44432
rect 71044 44368 71060 44432
rect 71124 44368 71140 44432
rect 71204 44368 71220 44432
rect 71284 44368 71322 44432
rect 70702 44352 71322 44368
rect 70702 44288 70740 44352
rect 70804 44288 70820 44352
rect 70884 44288 70900 44352
rect 70964 44288 70980 44352
rect 71044 44288 71060 44352
rect 71124 44288 71140 44352
rect 71204 44288 71220 44352
rect 71284 44288 71322 44352
rect 70702 34592 71322 44288
rect 70702 34528 70740 34592
rect 70804 34528 70820 34592
rect 70884 34528 70900 34592
rect 70964 34528 70980 34592
rect 71044 34528 71060 34592
rect 71124 34528 71140 34592
rect 71204 34528 71220 34592
rect 71284 34528 71322 34592
rect 70702 34512 71322 34528
rect 70702 34448 70740 34512
rect 70804 34448 70820 34512
rect 70884 34448 70900 34512
rect 70964 34448 70980 34512
rect 71044 34448 71060 34512
rect 71124 34448 71140 34512
rect 71204 34448 71220 34512
rect 71284 34448 71322 34512
rect 70702 34432 71322 34448
rect 70702 34368 70740 34432
rect 70804 34368 70820 34432
rect 70884 34368 70900 34432
rect 70964 34368 70980 34432
rect 71044 34368 71060 34432
rect 71124 34368 71140 34432
rect 71204 34368 71220 34432
rect 71284 34368 71322 34432
rect 70702 34352 71322 34368
rect 70702 34288 70740 34352
rect 70804 34288 70820 34352
rect 70884 34288 70900 34352
rect 70964 34288 70980 34352
rect 71044 34288 71060 34352
rect 71124 34288 71140 34352
rect 71204 34288 71220 34352
rect 71284 34288 71322 34352
rect 70702 24592 71322 34288
rect 70702 24528 70740 24592
rect 70804 24528 70820 24592
rect 70884 24528 70900 24592
rect 70964 24528 70980 24592
rect 71044 24528 71060 24592
rect 71124 24528 71140 24592
rect 71204 24528 71220 24592
rect 71284 24528 71322 24592
rect 70702 24512 71322 24528
rect 70702 24448 70740 24512
rect 70804 24448 70820 24512
rect 70884 24448 70900 24512
rect 70964 24448 70980 24512
rect 71044 24448 71060 24512
rect 71124 24448 71140 24512
rect 71204 24448 71220 24512
rect 71284 24448 71322 24512
rect 70702 24432 71322 24448
rect 70702 24368 70740 24432
rect 70804 24368 70820 24432
rect 70884 24368 70900 24432
rect 70964 24368 70980 24432
rect 71044 24368 71060 24432
rect 71124 24368 71140 24432
rect 71204 24368 71220 24432
rect 71284 24368 71322 24432
rect 70702 24352 71322 24368
rect 70702 24288 70740 24352
rect 70804 24288 70820 24352
rect 70884 24288 70900 24352
rect 70964 24288 70980 24352
rect 71044 24288 71060 24352
rect 71124 24288 71140 24352
rect 71204 24288 71220 24352
rect 71284 24288 71322 24352
rect 70702 14592 71322 24288
rect 70702 14528 70740 14592
rect 70804 14528 70820 14592
rect 70884 14528 70900 14592
rect 70964 14528 70980 14592
rect 71044 14528 71060 14592
rect 71124 14528 71140 14592
rect 71204 14528 71220 14592
rect 71284 14528 71322 14592
rect 70702 14512 71322 14528
rect 70702 14448 70740 14512
rect 70804 14448 70820 14512
rect 70884 14448 70900 14512
rect 70964 14448 70980 14512
rect 71044 14448 71060 14512
rect 71124 14448 71140 14512
rect 71204 14448 71220 14512
rect 71284 14448 71322 14512
rect 70702 14432 71322 14448
rect 70702 14368 70740 14432
rect 70804 14368 70820 14432
rect 70884 14368 70900 14432
rect 70964 14368 70980 14432
rect 71044 14368 71060 14432
rect 71124 14368 71140 14432
rect 71204 14368 71220 14432
rect 71284 14368 71322 14432
rect 70702 14352 71322 14368
rect 70702 14288 70740 14352
rect 70804 14288 70820 14352
rect 70884 14288 70900 14352
rect 70964 14288 70980 14352
rect 71044 14288 71060 14352
rect 71124 14288 71140 14352
rect 71204 14288 71220 14352
rect 71284 14288 71322 14352
rect 70702 4592 71322 14288
rect 70702 4528 70740 4592
rect 70804 4528 70820 4592
rect 70884 4528 70900 4592
rect 70964 4528 70980 4592
rect 71044 4528 71060 4592
rect 71124 4528 71140 4592
rect 71204 4528 71220 4592
rect 71284 4528 71322 4592
rect 70702 4512 71322 4528
rect 70702 4448 70740 4512
rect 70804 4448 70820 4512
rect 70884 4448 70900 4512
rect 70964 4448 70980 4512
rect 71044 4448 71060 4512
rect 71124 4448 71140 4512
rect 71204 4448 71220 4512
rect 71284 4448 71322 4512
rect 70702 4432 71322 4448
rect 70702 4368 70740 4432
rect 70804 4368 70820 4432
rect 70884 4368 70900 4432
rect 70964 4368 70980 4432
rect 71044 4368 71060 4432
rect 71124 4368 71140 4432
rect 71204 4368 71220 4432
rect 71284 4368 71322 4432
rect 70702 4352 71322 4368
rect 70702 4288 70740 4352
rect 70804 4288 70820 4352
rect 70884 4288 70900 4352
rect 70964 4288 70980 4352
rect 71044 4288 71060 4352
rect 71124 4288 71140 4352
rect 71204 4288 71220 4352
rect 71284 4288 71322 4352
rect 69059 3772 69125 3773
rect 69059 3708 69060 3772
rect 69124 3708 69125 3772
rect 69059 3707 69125 3708
rect 67702 2176 67740 2240
rect 67804 2176 67820 2240
rect 67884 2176 67900 2240
rect 67964 2176 67980 2240
rect 68044 2176 68060 2240
rect 68124 2176 68140 2240
rect 68204 2176 68220 2240
rect 68284 2176 68322 2240
rect 67702 2160 68322 2176
rect 67702 2096 67740 2160
rect 67804 2096 67820 2160
rect 67884 2096 67900 2160
rect 67964 2096 67980 2160
rect 68044 2096 68060 2160
rect 68124 2096 68140 2160
rect 68204 2096 68220 2160
rect 68284 2096 68322 2160
rect 67702 2080 68322 2096
rect 67702 2016 67740 2080
rect 67804 2016 67820 2080
rect 67884 2016 67900 2080
rect 67964 2016 67980 2080
rect 68044 2016 68060 2080
rect 68124 2016 68140 2080
rect 68204 2016 68220 2080
rect 68284 2016 68322 2080
rect 67702 2000 68322 2016
rect 67702 1936 67740 2000
rect 67804 1936 67820 2000
rect 67884 1936 67900 2000
rect 67964 1936 67980 2000
rect 68044 1936 68060 2000
rect 68124 1936 68140 2000
rect 68204 1936 68220 2000
rect 68284 1936 68322 2000
rect 65563 1324 65629 1325
rect 65563 1260 65564 1324
rect 65628 1260 65629 1324
rect 65563 1259 65629 1260
rect 67702 0 68322 1936
rect 70702 0 71322 4288
rect 73702 82240 74322 87000
rect 73702 82176 73740 82240
rect 73804 82176 73820 82240
rect 73884 82176 73900 82240
rect 73964 82176 73980 82240
rect 74044 82176 74060 82240
rect 74124 82176 74140 82240
rect 74204 82176 74220 82240
rect 74284 82176 74322 82240
rect 73702 82160 74322 82176
rect 73702 82096 73740 82160
rect 73804 82096 73820 82160
rect 73884 82096 73900 82160
rect 73964 82096 73980 82160
rect 74044 82096 74060 82160
rect 74124 82096 74140 82160
rect 74204 82096 74220 82160
rect 74284 82096 74322 82160
rect 73702 82080 74322 82096
rect 73702 82016 73740 82080
rect 73804 82016 73820 82080
rect 73884 82016 73900 82080
rect 73964 82016 73980 82080
rect 74044 82016 74060 82080
rect 74124 82016 74140 82080
rect 74204 82016 74220 82080
rect 74284 82016 74322 82080
rect 73702 82000 74322 82016
rect 73702 81936 73740 82000
rect 73804 81936 73820 82000
rect 73884 81936 73900 82000
rect 73964 81936 73980 82000
rect 74044 81936 74060 82000
rect 74124 81936 74140 82000
rect 74204 81936 74220 82000
rect 74284 81936 74322 82000
rect 73702 72240 74322 81936
rect 73702 72176 73740 72240
rect 73804 72176 73820 72240
rect 73884 72176 73900 72240
rect 73964 72176 73980 72240
rect 74044 72176 74060 72240
rect 74124 72176 74140 72240
rect 74204 72176 74220 72240
rect 74284 72176 74322 72240
rect 73702 72160 74322 72176
rect 73702 72096 73740 72160
rect 73804 72096 73820 72160
rect 73884 72096 73900 72160
rect 73964 72096 73980 72160
rect 74044 72096 74060 72160
rect 74124 72096 74140 72160
rect 74204 72096 74220 72160
rect 74284 72096 74322 72160
rect 73702 72080 74322 72096
rect 73702 72016 73740 72080
rect 73804 72016 73820 72080
rect 73884 72016 73900 72080
rect 73964 72016 73980 72080
rect 74044 72016 74060 72080
rect 74124 72016 74140 72080
rect 74204 72016 74220 72080
rect 74284 72016 74322 72080
rect 73702 72000 74322 72016
rect 73702 71936 73740 72000
rect 73804 71936 73820 72000
rect 73884 71936 73900 72000
rect 73964 71936 73980 72000
rect 74044 71936 74060 72000
rect 74124 71936 74140 72000
rect 74204 71936 74220 72000
rect 74284 71936 74322 72000
rect 73702 62240 74322 71936
rect 73702 62176 73740 62240
rect 73804 62176 73820 62240
rect 73884 62176 73900 62240
rect 73964 62176 73980 62240
rect 74044 62176 74060 62240
rect 74124 62176 74140 62240
rect 74204 62176 74220 62240
rect 74284 62176 74322 62240
rect 73702 62160 74322 62176
rect 73702 62096 73740 62160
rect 73804 62096 73820 62160
rect 73884 62096 73900 62160
rect 73964 62096 73980 62160
rect 74044 62096 74060 62160
rect 74124 62096 74140 62160
rect 74204 62096 74220 62160
rect 74284 62096 74322 62160
rect 73702 62080 74322 62096
rect 73702 62016 73740 62080
rect 73804 62016 73820 62080
rect 73884 62016 73900 62080
rect 73964 62016 73980 62080
rect 74044 62016 74060 62080
rect 74124 62016 74140 62080
rect 74204 62016 74220 62080
rect 74284 62016 74322 62080
rect 73702 62000 74322 62016
rect 73702 61936 73740 62000
rect 73804 61936 73820 62000
rect 73884 61936 73900 62000
rect 73964 61936 73980 62000
rect 74044 61936 74060 62000
rect 74124 61936 74140 62000
rect 74204 61936 74220 62000
rect 74284 61936 74322 62000
rect 73702 52240 74322 61936
rect 73702 52176 73740 52240
rect 73804 52176 73820 52240
rect 73884 52176 73900 52240
rect 73964 52176 73980 52240
rect 74044 52176 74060 52240
rect 74124 52176 74140 52240
rect 74204 52176 74220 52240
rect 74284 52176 74322 52240
rect 73702 52160 74322 52176
rect 73702 52096 73740 52160
rect 73804 52096 73820 52160
rect 73884 52096 73900 52160
rect 73964 52096 73980 52160
rect 74044 52096 74060 52160
rect 74124 52096 74140 52160
rect 74204 52096 74220 52160
rect 74284 52096 74322 52160
rect 73702 52080 74322 52096
rect 73702 52016 73740 52080
rect 73804 52016 73820 52080
rect 73884 52016 73900 52080
rect 73964 52016 73980 52080
rect 74044 52016 74060 52080
rect 74124 52016 74140 52080
rect 74204 52016 74220 52080
rect 74284 52016 74322 52080
rect 73702 52000 74322 52016
rect 73702 51936 73740 52000
rect 73804 51936 73820 52000
rect 73884 51936 73900 52000
rect 73964 51936 73980 52000
rect 74044 51936 74060 52000
rect 74124 51936 74140 52000
rect 74204 51936 74220 52000
rect 74284 51936 74322 52000
rect 73702 42240 74322 51936
rect 73702 42176 73740 42240
rect 73804 42176 73820 42240
rect 73884 42176 73900 42240
rect 73964 42176 73980 42240
rect 74044 42176 74060 42240
rect 74124 42176 74140 42240
rect 74204 42176 74220 42240
rect 74284 42176 74322 42240
rect 73702 42160 74322 42176
rect 73702 42096 73740 42160
rect 73804 42096 73820 42160
rect 73884 42096 73900 42160
rect 73964 42096 73980 42160
rect 74044 42096 74060 42160
rect 74124 42096 74140 42160
rect 74204 42096 74220 42160
rect 74284 42096 74322 42160
rect 73702 42080 74322 42096
rect 73702 42016 73740 42080
rect 73804 42016 73820 42080
rect 73884 42016 73900 42080
rect 73964 42016 73980 42080
rect 74044 42016 74060 42080
rect 74124 42016 74140 42080
rect 74204 42016 74220 42080
rect 74284 42016 74322 42080
rect 73702 42000 74322 42016
rect 73702 41936 73740 42000
rect 73804 41936 73820 42000
rect 73884 41936 73900 42000
rect 73964 41936 73980 42000
rect 74044 41936 74060 42000
rect 74124 41936 74140 42000
rect 74204 41936 74220 42000
rect 74284 41936 74322 42000
rect 73702 32240 74322 41936
rect 73702 32176 73740 32240
rect 73804 32176 73820 32240
rect 73884 32176 73900 32240
rect 73964 32176 73980 32240
rect 74044 32176 74060 32240
rect 74124 32176 74140 32240
rect 74204 32176 74220 32240
rect 74284 32176 74322 32240
rect 73702 32160 74322 32176
rect 73702 32096 73740 32160
rect 73804 32096 73820 32160
rect 73884 32096 73900 32160
rect 73964 32096 73980 32160
rect 74044 32096 74060 32160
rect 74124 32096 74140 32160
rect 74204 32096 74220 32160
rect 74284 32096 74322 32160
rect 73702 32080 74322 32096
rect 73702 32016 73740 32080
rect 73804 32016 73820 32080
rect 73884 32016 73900 32080
rect 73964 32016 73980 32080
rect 74044 32016 74060 32080
rect 74124 32016 74140 32080
rect 74204 32016 74220 32080
rect 74284 32016 74322 32080
rect 73702 32000 74322 32016
rect 73702 31936 73740 32000
rect 73804 31936 73820 32000
rect 73884 31936 73900 32000
rect 73964 31936 73980 32000
rect 74044 31936 74060 32000
rect 74124 31936 74140 32000
rect 74204 31936 74220 32000
rect 74284 31936 74322 32000
rect 73702 22240 74322 31936
rect 73702 22176 73740 22240
rect 73804 22176 73820 22240
rect 73884 22176 73900 22240
rect 73964 22176 73980 22240
rect 74044 22176 74060 22240
rect 74124 22176 74140 22240
rect 74204 22176 74220 22240
rect 74284 22176 74322 22240
rect 73702 22160 74322 22176
rect 73702 22096 73740 22160
rect 73804 22096 73820 22160
rect 73884 22096 73900 22160
rect 73964 22096 73980 22160
rect 74044 22096 74060 22160
rect 74124 22096 74140 22160
rect 74204 22096 74220 22160
rect 74284 22096 74322 22160
rect 73702 22080 74322 22096
rect 73702 22016 73740 22080
rect 73804 22016 73820 22080
rect 73884 22016 73900 22080
rect 73964 22016 73980 22080
rect 74044 22016 74060 22080
rect 74124 22016 74140 22080
rect 74204 22016 74220 22080
rect 74284 22016 74322 22080
rect 73702 22000 74322 22016
rect 73702 21936 73740 22000
rect 73804 21936 73820 22000
rect 73884 21936 73900 22000
rect 73964 21936 73980 22000
rect 74044 21936 74060 22000
rect 74124 21936 74140 22000
rect 74204 21936 74220 22000
rect 74284 21936 74322 22000
rect 73702 12240 74322 21936
rect 73702 12176 73740 12240
rect 73804 12176 73820 12240
rect 73884 12176 73900 12240
rect 73964 12176 73980 12240
rect 74044 12176 74060 12240
rect 74124 12176 74140 12240
rect 74204 12176 74220 12240
rect 74284 12176 74322 12240
rect 73702 12160 74322 12176
rect 73702 12096 73740 12160
rect 73804 12096 73820 12160
rect 73884 12096 73900 12160
rect 73964 12096 73980 12160
rect 74044 12096 74060 12160
rect 74124 12096 74140 12160
rect 74204 12096 74220 12160
rect 74284 12096 74322 12160
rect 73702 12080 74322 12096
rect 73702 12016 73740 12080
rect 73804 12016 73820 12080
rect 73884 12016 73900 12080
rect 73964 12016 73980 12080
rect 74044 12016 74060 12080
rect 74124 12016 74140 12080
rect 74204 12016 74220 12080
rect 74284 12016 74322 12080
rect 73702 12000 74322 12016
rect 73702 11936 73740 12000
rect 73804 11936 73820 12000
rect 73884 11936 73900 12000
rect 73964 11936 73980 12000
rect 74044 11936 74060 12000
rect 74124 11936 74140 12000
rect 74204 11936 74220 12000
rect 74284 11936 74322 12000
rect 73702 2240 74322 11936
rect 73702 2176 73740 2240
rect 73804 2176 73820 2240
rect 73884 2176 73900 2240
rect 73964 2176 73980 2240
rect 74044 2176 74060 2240
rect 74124 2176 74140 2240
rect 74204 2176 74220 2240
rect 74284 2176 74322 2240
rect 73702 2160 74322 2176
rect 73702 2096 73740 2160
rect 73804 2096 73820 2160
rect 73884 2096 73900 2160
rect 73964 2096 73980 2160
rect 74044 2096 74060 2160
rect 74124 2096 74140 2160
rect 74204 2096 74220 2160
rect 74284 2096 74322 2160
rect 73702 2080 74322 2096
rect 73702 2016 73740 2080
rect 73804 2016 73820 2080
rect 73884 2016 73900 2080
rect 73964 2016 73980 2080
rect 74044 2016 74060 2080
rect 74124 2016 74140 2080
rect 74204 2016 74220 2080
rect 74284 2016 74322 2080
rect 73702 2000 74322 2016
rect 73702 1936 73740 2000
rect 73804 1936 73820 2000
rect 73884 1936 73900 2000
rect 73964 1936 73980 2000
rect 74044 1936 74060 2000
rect 74124 1936 74140 2000
rect 74204 1936 74220 2000
rect 74284 1936 74322 2000
rect 73702 0 74322 1936
use sky130_fd_sc_hd__clkinv_4  _10_
timestamp 1
transform -1 0 43056 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _11_
timestamp 1
transform 1 0 28336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _12_
timestamp 1
transform -1 0 40848 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _13_
timestamp 1
transform 1 0 33580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _14_
timestamp 1
transform 1 0 32108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _15_
timestamp 1
transform 1 0 31740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _16_
timestamp 1
transform 1 0 31188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _17_
timestamp 1
transform 1 0 30912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _18_
timestamp 1
transform 1 0 31004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_2  _19_
timestamp 1
transform 1 0 30360 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_2  _20_
timestamp 1
transform 1 0 30176 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_2  _21_
timestamp 1
transform 1 0 29348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_2  _22_
timestamp 1
transform 1 0 29532 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _23_
timestamp 1
transform 1 0 46644 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _24_
timestamp 1
transform 1 0 48208 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _25_
timestamp 1
transform 1 0 49864 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _26_
timestamp 1
transform 1 0 51428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _27_
timestamp 1
transform 1 0 52900 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _28_
timestamp 1
transform 1 0 54556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _29_
timestamp 1
transform 1 0 56028 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _30_
timestamp 1
transform 1 0 57776 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _31_
timestamp 1
transform 1 0 59064 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _32_
timestamp 1
transform 1 0 60536 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _33_
timestamp 1
transform 1 0 62008 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _34_
timestamp 1
transform 1 0 63480 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _35_
timestamp 1
transform 1 0 64952 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _36_
timestamp 1
transform 1 0 66424 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _37_
timestamp 1
transform 1 0 68080 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _38_
timestamp 1
transform 1 0 69184 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _39_
timestamp 1
transform -1 0 35788 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _40_
timestamp 1
transform -1 0 35052 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _41_
timestamp 1
transform -1 0 35420 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _42_
timestamp 1
transform -1 0 34132 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _43_
timestamp 1
transform -1 0 35328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _44_
timestamp 1
transform 1 0 32844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _45_
timestamp 1
transform -1 0 35052 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform 1 0 35788 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform -1 0 35236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform -1 0 35236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 31096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform -1 0 33028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform -1 0 31188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform -1 0 30360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform 1 0 30360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform -1 0 30176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform -1 0 46644 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform -1 0 46828 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform -1 0 48208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform -1 0 49864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform -1 0 51428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform -1 0 35788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform -1 0 53084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform -1 0 54556 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1
transform -1 0 56028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1
transform -1 0 59248 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1
transform -1 0 59248 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1
transform -1 0 59248 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1
transform -1 0 59248 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1
transform -1 0 59248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1
transform -1 0 59248 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1
transform -1 0 59248 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1
transform 1 0 59616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1
transform -1 0 59248 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1
transform 1 0 59432 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1
transform 1 0 59248 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1
transform -1 0 60720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1
transform -1 0 60720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1
transform -1 0 60720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1
transform -1 0 60720 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1
transform -1 0 60720 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1
transform 1 0 61088 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1
transform -1 0 60720 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1
transform 1 0 60904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1
transform -1 0 60720 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1
transform 1 0 60720 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1
transform -1 0 60720 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1
transform -1 0 62192 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1
transform -1 0 62192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1
transform -1 0 62192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1
transform -1 0 62192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1
transform -1 0 62192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1
transform -1 0 62192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1
transform -1 0 62192 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1
transform 1 0 62560 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1
transform -1 0 62192 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1
transform 1 0 62376 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1
transform 1 0 62192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1
transform 1 0 63480 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1
transform 1 0 63480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1
transform 1 0 63480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1
transform 1 0 63480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1
transform 1 0 63480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_57
timestamp 1
transform 1 0 63480 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_58
timestamp 1
transform 1 0 63480 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_59
timestamp 1
transform 1 0 63848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_60
timestamp 1
transform -1 0 63664 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_61
timestamp 1
transform 1 0 63664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_62
timestamp 1
transform -1 0 65872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_63
timestamp 1
transform -1 0 65136 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_64
timestamp 1
transform 1 0 66424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_65
timestamp 1
transform 1 0 66424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_66
timestamp 1
transform 1 0 66424 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_67
timestamp 1
transform 1 0 66424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_68
timestamp 1
transform 1 0 66424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_69
timestamp 1
transform 1 0 66424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_70
timestamp 1
transform 1 0 66424 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_71
timestamp 1
transform 1 0 66424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_72
timestamp 1
transform -1 0 66608 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_73
timestamp 1
transform 1 0 66424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_74
timestamp 1
transform 1 0 66424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_75
timestamp 1
transform 1 0 35420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_76
timestamp 1
transform -1 0 68264 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_77
timestamp 1
transform 1 0 69184 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_78
timestamp 1
transform 1 0 69184 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_79
timestamp 1
transform 1 0 69184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_80
timestamp 1
transform 1 0 69184 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_81
timestamp 1
transform 1 0 69184 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_82
timestamp 1
transform 1 0 69184 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_83
timestamp 1
transform 1 0 69184 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_84
timestamp 1
transform 1 0 69184 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_85
timestamp 1
transform -1 0 69368 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_86
timestamp 1
transform 1 0 69184 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_87
timestamp 1
transform 1 0 69184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_88
timestamp 1
transform -1 0 32844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_89
timestamp 1
transform -1 0 34776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_90
timestamp 1
transform 1 0 36524 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_91
timestamp 1
transform -1 0 33212 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_92
timestamp 1
transform -1 0 32292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_93
timestamp 1
transform 1 0 32476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_94
timestamp 1
transform -1 0 31924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_95
timestamp 1
transform -1 0 31372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_96
timestamp 1
transform 1 0 65688 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_97
timestamp 1
transform -1 0 44068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_98
timestamp 1
transform -1 0 48392 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_99
timestamp 1
transform -1 0 48944 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_100
timestamp 1
transform -1 0 34316 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_101
timestamp 1
transform -1 0 34500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_102
timestamp 1
transform -1 0 33028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_103
timestamp 1
transform -1 0 65872 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_104
timestamp 1
transform -1 0 66056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_105
timestamp 1
transform -1 0 65872 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_106
timestamp 1
transform 1 0 44620 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1
transform 1 0 65688 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1
transform -1 0 47380 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1
transform 1 0 65688 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_16  clkload0
timestamp 1
transform -1 0 47380 0 1 5440
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_2  fanout84
timestamp 1
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout85
timestamp 1
transform -1 0 32568 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout86
timestamp 1
transform -1 0 30912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout87
timestamp 1
transform 1 0 30268 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout88
timestamp 1
transform -1 0 30268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout89
timestamp 1
transform -1 0 31648 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_3
timestamp 1562078211
transform 1 0 1288 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_15
timestamp 1562078211
transform 1 0 2392 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3496 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_29
timestamp 1562078211
transform 1 0 3680 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_41
timestamp 1562078211
transform 1 0 4784 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1
transform 1 0 5888 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1
transform 1 0 6072 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_57
timestamp 1562078211
transform 1 0 6256 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_69
timestamp 1562078211
transform 1 0 7360 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_81
timestamp 1
transform 1 0 8464 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1
transform 1 0 8648 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_85
timestamp 1562078211
transform 1 0 8832 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_97
timestamp 1562078211
transform 1 0 9936 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109
timestamp 1
transform 1 0 11040 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1
transform 1 0 11224 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_113
timestamp 1562078211
transform 1 0 11408 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_125
timestamp 1562078211
transform 1 0 12512 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1
transform 1 0 13616 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1
transform 1 0 13800 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_141
timestamp 1562078211
transform 1 0 13984 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_153
timestamp 1562078211
transform 1 0 15088 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1
transform 1 0 16192 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1
transform 1 0 16376 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_169
timestamp 1562078211
transform 1 0 16560 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_181
timestamp 1562078211
transform 1 0 17664 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1
transform 1 0 18768 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1
transform 1 0 18952 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_197
timestamp 1562078211
transform 1 0 19136 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_209
timestamp 1562078211
transform 1 0 20240 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1
transform 1 0 21344 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1
transform 1 0 21528 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_225
timestamp 1562078211
transform 1 0 21712 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_0_237
timestamp 1
transform 1 0 22816 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_248
timestamp 1
transform 1 0 23828 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_269
timestamp 1
transform 1 0 25760 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_271
timestamp 1
transform 1 0 25944 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1
transform 1 0 26864 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_283
timestamp 1
transform 1 0 27048 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1
transform 1 0 29440 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_311
timestamp 1
transform 1 0 29624 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_361
timestamp 1
transform 1 0 34224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1
transform 1 0 34408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1
transform 1 0 34592 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1
transform 1 0 36984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1
transform 1 0 37168 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_395
timestamp 1
transform 1 0 37352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_445
timestamp 1
transform 1 0 41952 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1
transform 1 0 42136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_473
timestamp 1
transform 1 0 44528 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1
transform 1 0 44712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1
transform 1 0 44896 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_479
timestamp 1
transform 1 0 45080 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_529
timestamp 1
transform 1 0 49680 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1
transform 1 0 49864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_557
timestamp 1
transform 1 0 52256 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1
transform 1 0 52440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_585
timestamp 1
transform 1 0 54832 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1
transform 1 0 55016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_613
timestamp 1
transform 1 0 57408 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1
transform 1 0 57592 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_0_617
timestamp 1562078211
transform 1 0 57776 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_629
timestamp 1
transform 1 0 58880 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_641
timestamp 1
transform 1 0 59984 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_643
timestamp 1
transform 1 0 60168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_645
timestamp 1
transform 1 0 60352 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_649
timestamp 1
transform 1 0 60720 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_653
timestamp 1
transform 1 0 61088 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_665
timestamp 1
transform 1 0 62192 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_669
timestamp 1
transform 1 0 62560 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 1
transform 1 0 62744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_0_673
timestamp 1
transform 1 0 62928 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_677
timestamp 1
transform 1 0 63296 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_697
timestamp 1
transform 1 0 65136 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1
transform 1 0 65320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_709
timestamp 1
transform 1 0 66240 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_713
timestamp 1
transform 1 0 66608 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_725
timestamp 1
transform 1 0 67712 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_727
timestamp 1
transform 1 0 67896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_0_735
timestamp 1
transform 1 0 68632 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_739
timestamp 1
transform 1 0 69000 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_743
timestamp 1
transform 1 0 69368 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_753
timestamp 1
transform 1 0 70288 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 1
transform 1 0 70472 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_781
timestamp 1
transform 1 0 72864 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_783
timestamp 1
transform 1 0 73048 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_0_793
timestamp 1
transform 1 0 73968 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_3
timestamp 1562078211
transform 1 0 1288 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_15
timestamp 1562078211
transform 1 0 2392 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_27
timestamp 1562078211
transform 1 0 3496 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_39
timestamp 1562078211
transform 1 0 4600 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_51
timestamp 1
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6072 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_57
timestamp 1562078211
transform 1 0 6256 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_69
timestamp 1562078211
transform 1 0 7360 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_81
timestamp 1562078211
transform 1 0 8464 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_93
timestamp 1562078211
transform 1 0 9568 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_105
timestamp 1
transform 1 0 10672 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_109
timestamp 1
transform 1 0 11040 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11224 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_113
timestamp 1562078211
transform 1 0 11408 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_125
timestamp 1562078211
transform 1 0 12512 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_137
timestamp 1562078211
transform 1 0 13616 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_149
timestamp 1562078211
transform 1 0 14720 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_161
timestamp 1
transform 1 0 15824 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_165
timestamp 1
transform 1 0 16192 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16376 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_169
timestamp 1562078211
transform 1 0 16560 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_181
timestamp 1562078211
transform 1 0 17664 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_193
timestamp 1562078211
transform 1 0 18768 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_205
timestamp 1562078211
transform 1 0 19872 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_217
timestamp 1
transform 1 0 20976 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1
transform 1 0 21344 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21528 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_225
timestamp 1562078211
transform 1 0 21712 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_237
timestamp 1562078211
transform 1 0 22816 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1
transform 1 0 23920 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_251
timestamp 1
transform 1 0 24104 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_301
timestamp 1
transform 1 0 28704 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_303
timestamp 1
transform 1 0 28888 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1
transform 1 0 32016 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_339
timestamp 1
transform 1 0 32200 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_356
timestamp 1
transform 1 0 33764 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1
transform 1 0 42136 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_449
timestamp 1
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_490
timestamp 1
transform 1 0 46092 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_509
timestamp 1
transform 1 0 47840 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_556
timestamp 1
transform 1 0 52164 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_569
timestamp 1
transform 1 0 53360 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_625
timestamp 1
transform 1 0 58512 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_629
timestamp 1
transform 1 0 58880 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_633
timestamp 1
transform 1 0 59248 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_643
timestamp 1
transform 1 0 60168 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_657
timestamp 1
transform 1 0 61456 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_661
timestamp 1
transform 1 0 61824 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1
transform 1 0 62744 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_673
timestamp 1
transform 1 0 62928 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_677
timestamp 1
transform 1 0 63296 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_697
timestamp 1
transform 1 0 65136 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_701
timestamp 1
transform 1 0 65504 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1
transform 1 0 67896 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_729
timestamp 1
transform 1 0 68080 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_781
timestamp 1
transform 1 0 72864 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1
transform 1 0 73048 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_1_785
timestamp 1562078211
transform 1 0 73232 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_1_797
timestamp 1
transform 1 0 74336 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_3
timestamp 1562078211
transform 1 0 1288 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_15
timestamp 1562078211
transform 1 0 2392 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3496 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_29
timestamp 1562078211
transform 1 0 3680 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_41
timestamp 1562078211
transform 1 0 4784 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_53
timestamp 1562078211
transform 1 0 5888 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_65
timestamp 1562078211
transform 1 0 6992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_77
timestamp 1
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8648 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_85
timestamp 1562078211
transform 1 0 8832 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_97
timestamp 1562078211
transform 1 0 9936 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_109
timestamp 1562078211
transform 1 0 11040 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_121
timestamp 1562078211
transform 1 0 12144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_133
timestamp 1
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_137
timestamp 1
transform 1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13800 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_141
timestamp 1562078211
transform 1 0 13984 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_153
timestamp 1562078211
transform 1 0 15088 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_165
timestamp 1562078211
transform 1 0 16192 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_177
timestamp 1562078211
transform 1 0 17296 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_189
timestamp 1
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_193
timestamp 1
transform 1 0 18768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 18952 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_197
timestamp 1562078211
transform 1 0 19136 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_209
timestamp 1562078211
transform 1 0 20240 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_221
timestamp 1562078211
transform 1 0 21344 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_233
timestamp 1562078211
transform 1 0 22448 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_2_245
timestamp 1
transform 1 0 23552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_249
timestamp 1
transform 1 0 23920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24104 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_253
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_257
timestamp 1
transform 1 0 24656 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_259
timestamp 1
transform 1 0 24840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_296
timestamp 1
transform 1 0 28244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1
transform 1 0 34408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_365
timestamp 1
transform 1 0 34592 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_369
timestamp 1
transform 1 0 34960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_378
timestamp 1
transform 1 0 35788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_388
timestamp 1
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_408
timestamp 1
transform 1 0 38548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1
transform 1 0 39468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_421
timestamp 1
transform 1 0 39744 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_431
timestamp 1
transform 1 0 40664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_433
timestamp 1
transform 1 0 40848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1
transform 1 0 44620 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1
transform 1 0 44896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_491
timestamp 1
transform 1 0 46184 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_501
timestamp 1
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_513
timestamp 1
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_529
timestamp 1
transform 1 0 49680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1
transform 1 0 49864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_533
timestamp 1
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_2_542
timestamp 1
transform 1 0 50876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_2_564
timestamp 1
transform 1 0 52900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_568
timestamp 1
transform 1 0 53268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_570
timestamp 1
transform 1 0 53452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_585
timestamp 1
transform 1 0 54832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1
transform 1 0 55016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_597
timestamp 1
transform 1 0 55936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_599
timestamp 1
transform 1 0 56120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_614
timestamp 1
transform 1 0 57500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_641
timestamp 1
transform 1 0 59984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1
transform 1 0 60168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_645
timestamp 1
transform 1 0 60352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_673
timestamp 1
transform 1 0 62928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_677
timestamp 1
transform 1 0 63296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_697
timestamp 1
transform 1 0 65136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1
transform 1 0 65320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_709
timestamp 1
transform 1 0 66240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_735
timestamp 1
transform 1 0 68632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_739
timestamp 1
transform 1 0 69000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_751
timestamp 1
transform 1 0 70104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1
transform 1 0 70472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_771
timestamp 1
transform 1 0 71944 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_2_779
timestamp 1562078211
transform 1 0 72680 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_2_791
timestamp 1
transform 1 0 73784 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_799
timestamp 1
transform 1 0 74520 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_3
timestamp 1562078211
transform 1 0 1288 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_15
timestamp 1562078211
transform 1 0 2392 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_27
timestamp 1562078211
transform 1 0 3496 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_39
timestamp 1562078211
transform 1 0 4600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_51
timestamp 1
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6072 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_57
timestamp 1562078211
transform 1 0 6256 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_69
timestamp 1562078211
transform 1 0 7360 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_81
timestamp 1562078211
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_93
timestamp 1562078211
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_105
timestamp 1
transform 1 0 10672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1
transform 1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11224 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_113
timestamp 1562078211
transform 1 0 11408 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_125
timestamp 1562078211
transform 1 0 12512 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_137
timestamp 1562078211
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_149
timestamp 1562078211
transform 1 0 14720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_161
timestamp 1
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1
transform 1 0 16192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16376 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_169
timestamp 1562078211
transform 1 0 16560 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_181
timestamp 1562078211
transform 1 0 17664 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_193
timestamp 1562078211
transform 1 0 18768 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_205
timestamp 1562078211
transform 1 0 19872 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_217
timestamp 1
transform 1 0 20976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1
transform 1 0 21344 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21528 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_225
timestamp 1562078211
transform 1 0 21712 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_237
timestamp 1562078211
transform 1 0 22816 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_249
timestamp 1562078211
transform 1 0 23920 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_261
timestamp 1
transform 1 0 25024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_265
timestamp 1
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_267
timestamp 1
transform 1 0 25576 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_281
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_285
timestamp 1
transform 1 0 27232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_330
timestamp 1
transform 1 0 31372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_337
timestamp 1
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_372
timestamp 1
transform 1 0 35236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_388
timestamp 1
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_407
timestamp 1
transform 1 0 38456 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_415
timestamp 1562078211
transform 1 0 39192 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_3_427
timestamp 1
transform 1 0 40296 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_435
timestamp 1
transform 1 0 41032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_457
timestamp 1
transform 1 0 43056 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_465
timestamp 1
transform 1 0 43792 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_484
timestamp 1562078211
transform 1 0 45540 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_3_496
timestamp 1
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_505
timestamp 1562078211
transform 1 0 47472 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_517
timestamp 1562078211
transform 1 0 48576 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_529
timestamp 1562078211
transform 1 0 49680 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_541
timestamp 1562078211
transform 1 0 50784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_553
timestamp 1
transform 1 0 51888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_557
timestamp 1
transform 1 0 52256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1
transform 1 0 52440 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_561
timestamp 1562078211
transform 1 0 52624 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_573
timestamp 1562078211
transform 1 0 53728 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_585
timestamp 1562078211
transform 1 0 54832 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_597
timestamp 1562078211
transform 1 0 55936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_609
timestamp 1
transform 1 0 57040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_613
timestamp 1
transform 1 0 57408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1
transform 1 0 57592 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_623
timestamp 1
transform 1 0 58328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_639
timestamp 1
transform 1 0 59800 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_649
timestamp 1562078211
transform 1 0 60720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_661
timestamp 1
transform 1 0 61824 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_665
timestamp 1
transform 1 0 62192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_669
timestamp 1
transform 1 0 62560 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1
transform 1 0 62744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_673
timestamp 1
transform 1 0 62928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_677
timestamp 1
transform 1 0 63296 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_681
timestamp 1
transform 1 0 63664 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_707
timestamp 1
transform 1 0 66056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_713
timestamp 1
transform 1 0 66608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_717
timestamp 1
transform 1 0 66976 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_726
timestamp 1
transform 1 0 67804 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_729
timestamp 1562078211
transform 1 0 68080 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_759
timestamp 1562078211
transform 1 0 70840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_771
timestamp 1562078211
transform 1 0 71944 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1
transform 1 0 73048 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_3_785
timestamp 1562078211
transform 1 0 73232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_3_797
timestamp 1
transform 1 0 74336 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_3
timestamp 1562078211
transform 1 0 1288 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_15
timestamp 1562078211
transform 1 0 2392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3496 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_29
timestamp 1562078211
transform 1 0 3680 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_41
timestamp 1562078211
transform 1 0 4784 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_53
timestamp 1562078211
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_65
timestamp 1562078211
transform 1 0 6992 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_77
timestamp 1
transform 1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1
transform 1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8648 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_85
timestamp 1562078211
transform 1 0 8832 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_97
timestamp 1562078211
transform 1 0 9936 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_109
timestamp 1562078211
transform 1 0 11040 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_121
timestamp 1562078211
transform 1 0 12144 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_133
timestamp 1
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1
transform 1 0 13616 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13800 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_141
timestamp 1562078211
transform 1 0 13984 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_153
timestamp 1562078211
transform 1 0 15088 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_165
timestamp 1562078211
transform 1 0 16192 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_177
timestamp 1562078211
transform 1 0 17296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_189
timestamp 1
transform 1 0 18400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1
transform 1 0 18768 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 18952 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_197
timestamp 1562078211
transform 1 0 19136 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_209
timestamp 1562078211
transform 1 0 20240 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_221
timestamp 1562078211
transform 1 0 21344 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_233
timestamp 1562078211
transform 1 0 22448 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_245
timestamp 1
transform 1 0 23552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_249
timestamp 1
transform 1 0 23920 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24104 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_253
timestamp 1562078211
transform 1 0 24288 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_265
timestamp 1562078211
transform 1 0 25392 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_277
timestamp 1
transform 1 0 26496 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_365
timestamp 1
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_378
timestamp 1
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_391
timestamp 1
transform 1 0 36984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_395
timestamp 1
transform 1 0 37352 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_397
timestamp 1
transform 1 0 37536 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_404
timestamp 1562078211
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_416
timestamp 1
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_421
timestamp 1562078211
transform 1 0 39744 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_433
timestamp 1
transform 1 0 40848 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_443
timestamp 1562078211
transform 1 0 41768 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_455
timestamp 1562078211
transform 1 0 42872 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_4_467
timestamp 1
transform 1 0 43976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1
transform 1 0 44712 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_477
timestamp 1562078211
transform 1 0 44896 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_489
timestamp 1
transform 1 0 46000 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_493
timestamp 1
transform 1 0 46368 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_495
timestamp 1
transform 1 0 46552 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_498
timestamp 1562078211
transform 1 0 46828 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_510
timestamp 1562078211
transform 1 0 47932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_4_522
timestamp 1
transform 1 0 49036 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_530
timestamp 1
transform 1 0 49772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_533
timestamp 1562078211
transform 1 0 50048 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_545
timestamp 1562078211
transform 1 0 51152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_557
timestamp 1
transform 1 0 52256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_561
timestamp 1
transform 1 0 52624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_563
timestamp 1
transform 1 0 52808 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_566
timestamp 1562078211
transform 1 0 53084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_4_578
timestamp 1
transform 1 0 54188 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_586
timestamp 1
transform 1 0 54924 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_589
timestamp 1562078211
transform 1 0 55200 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_601
timestamp 1562078211
transform 1 0 56304 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_613
timestamp 1
transform 1 0 57408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_4_633
timestamp 1
transform 1 0 59248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_641
timestamp 1
transform 1 0 59984 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1
transform 1 0 60168 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_645
timestamp 1
transform 1 0 60352 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_649
timestamp 1562078211
transform 1 0 60720 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_661
timestamp 1
transform 1 0 61824 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_665
timestamp 1562078211
transform 1 0 62192 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_677
timestamp 1
transform 1 0 63296 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_689
timestamp 1
transform 1 0 64400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_693
timestamp 1
transform 1 0 64768 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_697
timestamp 1
transform 1 0 65136 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1
transform 1 0 65320 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_707
timestamp 1
transform 1 0 66056 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_713
timestamp 1562078211
transform 1 0 66608 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_4_725
timestamp 1
transform 1 0 67712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_4_731
timestamp 1
transform 1 0 68264 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_739
timestamp 1
transform 1 0 69000 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_743
timestamp 1562078211
transform 1 0 69368 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1
transform 1 0 70472 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_757
timestamp 1562078211
transform 1 0 70656 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_769
timestamp 1562078211
transform 1 0 71760 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_4_781
timestamp 1562078211
transform 1 0 72864 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_4_793
timestamp 1
transform 1 0 73968 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_3
timestamp 1562078211
transform 1 0 1288 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_15
timestamp 1562078211
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_27
timestamp 1562078211
transform 1 0 3496 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_39
timestamp 1562078211
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_51
timestamp 1
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6072 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_57
timestamp 1562078211
transform 1 0 6256 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_69
timestamp 1562078211
transform 1 0 7360 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_81
timestamp 1562078211
transform 1 0 8464 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_93
timestamp 1562078211
transform 1 0 9568 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_105
timestamp 1
transform 1 0 10672 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11224 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_113
timestamp 1562078211
transform 1 0 11408 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_125
timestamp 1562078211
transform 1 0 12512 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_137
timestamp 1562078211
transform 1 0 13616 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_149
timestamp 1562078211
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_161
timestamp 1
transform 1 0 15824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1
transform 1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16376 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_169
timestamp 1562078211
transform 1 0 16560 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_181
timestamp 1562078211
transform 1 0 17664 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_193
timestamp 1562078211
transform 1 0 18768 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_205
timestamp 1562078211
transform 1 0 19872 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_217
timestamp 1
transform 1 0 20976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21528 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_225
timestamp 1562078211
transform 1 0 21712 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_237
timestamp 1562078211
transform 1 0 22816 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_249
timestamp 1562078211
transform 1 0 23920 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_261
timestamp 1562078211
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_273
timestamp 1
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_277
timestamp 1
transform 1 0 26496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_281
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_285
timestamp 1
transform 1 0 27232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_287
timestamp 1
transform 1 0 27416 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_296
timestamp 1
transform 1 0 28244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_337
timestamp 1
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_348
timestamp 1
transform 1 0 33028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_388
timestamp 1
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_393
timestamp 1562078211
transform 1 0 37168 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_405
timestamp 1562078211
transform 1 0 38272 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_5_417
timestamp 1
transform 1 0 39376 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_425
timestamp 1
transform 1 0 40112 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_433
timestamp 1562078211
transform 1 0 40848 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_445
timestamp 1
transform 1 0 41952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1
transform 1 0 42136 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_449
timestamp 1562078211
transform 1 0 42320 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_461
timestamp 1562078211
transform 1 0 43424 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_473
timestamp 1562078211
transform 1 0 44528 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_5_485
timestamp 1
transform 1 0 45632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_493
timestamp 1
transform 1 0 46368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_505
timestamp 1
transform 1 0 47472 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_509
timestamp 1
transform 1 0 47840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_5_521
timestamp 1
transform 1 0 48944 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_539
timestamp 1
transform 1 0 50600 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_543
timestamp 1
transform 1 0 50968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_545
timestamp 1
transform 1 0 51152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_556
timestamp 1
transform 1 0 52164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_561
timestamp 1
transform 1 0 52624 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_563
timestamp 1
transform 1 0 52808 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_572
timestamp 1
transform 1 0 53636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_590
timestamp 1
transform 1 0 55292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_594
timestamp 1
transform 1 0 55660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_5_606
timestamp 1
transform 1 0 56764 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_614
timestamp 1
transform 1 0 57500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_5_625
timestamp 1
transform 1 0 58512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_629
timestamp 1
transform 1 0 58880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_5_639
timestamp 1
transform 1 0 59800 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_649
timestamp 1562078211
transform 1 0 60720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_661
timestamp 1
transform 1 0 61824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1
transform 1 0 62744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_673
timestamp 1
transform 1 0 62928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_677
timestamp 1
transform 1 0 63296 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_5_687
timestamp 1
transform 1 0 64216 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_703
timestamp 1
transform 1 0 65688 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_719
timestamp 1
transform 1 0 67160 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1
transform 1 0 67896 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_737
timestamp 1
transform 1 0 68816 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_749
timestamp 1562078211
transform 1 0 69920 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_761
timestamp 1562078211
transform 1 0 71024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_5_773
timestamp 1
transform 1 0 72128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_781
timestamp 1
transform 1 0 72864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1
transform 1 0 73048 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_5_785
timestamp 1562078211
transform 1 0 73232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_5_797
timestamp 1
transform 1 0 74336 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_3
timestamp 1562078211
transform 1 0 1288 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_15
timestamp 1562078211
transform 1 0 2392 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3496 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_29
timestamp 1562078211
transform 1 0 3680 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_41
timestamp 1562078211
transform 1 0 4784 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_53
timestamp 1562078211
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_65
timestamp 1562078211
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_77
timestamp 1
transform 1 0 8096 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8648 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_85
timestamp 1562078211
transform 1 0 8832 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_97
timestamp 1562078211
transform 1 0 9936 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_109
timestamp 1562078211
transform 1 0 11040 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_121
timestamp 1562078211
transform 1 0 12144 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_133
timestamp 1
transform 1 0 13248 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1
transform 1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13800 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_141
timestamp 1562078211
transform 1 0 13984 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_153
timestamp 1562078211
transform 1 0 15088 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_165
timestamp 1562078211
transform 1 0 16192 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_177
timestamp 1562078211
transform 1 0 17296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_189
timestamp 1
transform 1 0 18400 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1
transform 1 0 18768 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 18952 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_197
timestamp 1562078211
transform 1 0 19136 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_209
timestamp 1562078211
transform 1 0 20240 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_221
timestamp 1562078211
transform 1 0 21344 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_233
timestamp 1562078211
transform 1 0 22448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_245
timestamp 1
transform 1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_249
timestamp 1
transform 1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24104 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_253
timestamp 1562078211
transform 1 0 24288 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_265
timestamp 1562078211
transform 1 0 25392 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_277
timestamp 1562078211
transform 1 0 26496 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_6_289
timestamp 1
transform 1 0 27600 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_297
timestamp 1
transform 1 0 28336 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_309
timestamp 1
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_6_333
timestamp 1
transform 1 0 31648 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_337
timestamp 1
transform 1 0 32016 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_346
timestamp 1
transform 1 0 32844 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_354
timestamp 1
transform 1 0 33580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1
transform 1 0 34316 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_379
timestamp 1562078211
transform 1 0 35880 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_391
timestamp 1562078211
transform 1 0 36984 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_403
timestamp 1562078211
transform 1 0 38088 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_415
timestamp 1
transform 1 0 39192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1
transform 1 0 39560 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_421
timestamp 1562078211
transform 1 0 39744 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_433
timestamp 1562078211
transform 1 0 40848 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_445
timestamp 1562078211
transform 1 0 41952 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_457
timestamp 1562078211
transform 1 0 43056 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_469
timestamp 1
transform 1 0 44160 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_473
timestamp 1
transform 1 0 44528 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1
transform 1 0 44712 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_6_477
timestamp 1
transform 1 0 44896 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_481
timestamp 1
transform 1 0 45264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_483
timestamp 1
transform 1 0 45448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_6_500
timestamp 1
transform 1 0 47012 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_504
timestamp 1
transform 1 0 47380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_521
timestamp 1
transform 1 0 48944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_529
timestamp 1
transform 1 0 49680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1
transform 1 0 49864 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_533
timestamp 1562078211
transform 1 0 50048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_545
timestamp 1562078211
transform 1 0 51152 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_557
timestamp 1562078211
transform 1 0 52256 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_569
timestamp 1562078211
transform 1 0 53360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_581
timestamp 1
transform 1 0 54464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_585
timestamp 1
transform 1 0 54832 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1
transform 1 0 55016 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_589
timestamp 1562078211
transform 1 0 55200 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_601
timestamp 1562078211
transform 1 0 56304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_613
timestamp 1562078211
transform 1 0 57408 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_625
timestamp 1
transform 1 0 58512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_629
timestamp 1
transform 1 0 58880 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_6_633
timestamp 1
transform 1 0 59248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_641
timestamp 1
transform 1 0 59984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1
transform 1 0 60168 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_645
timestamp 1
transform 1 0 60352 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_6_655
timestamp 1
transform 1 0 61272 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_665
timestamp 1562078211
transform 1 0 62192 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_677
timestamp 1
transform 1 0 63296 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_681
timestamp 1562078211
transform 1 0 63664 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_693
timestamp 1
transform 1 0 64768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_697
timestamp 1
transform 1 0 65136 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1
transform 1 0 65320 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_701
timestamp 1
transform 1 0 65504 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_709
timestamp 1
transform 1 0 66240 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_713
timestamp 1562078211
transform 1 0 66608 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_725
timestamp 1562078211
transform 1 0 67712 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_6_737
timestamp 1
transform 1 0 68816 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_743
timestamp 1562078211
transform 1 0 69368 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1
transform 1 0 70472 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_757
timestamp 1562078211
transform 1 0 70656 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_769
timestamp 1562078211
transform 1 0 71760 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_6_781
timestamp 1562078211
transform 1 0 72864 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_6_793
timestamp 1
transform 1 0 73968 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_3
timestamp 1562078211
transform 1 0 1288 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_15
timestamp 1562078211
transform 1 0 2392 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_27
timestamp 1562078211
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_39
timestamp 1562078211
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_51
timestamp 1
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6072 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_57
timestamp 1562078211
transform 1 0 6256 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_69
timestamp 1562078211
transform 1 0 7360 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_81
timestamp 1562078211
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_93
timestamp 1562078211
transform 1 0 9568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_105
timestamp 1
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11224 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_113
timestamp 1562078211
transform 1 0 11408 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_125
timestamp 1562078211
transform 1 0 12512 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_137
timestamp 1562078211
transform 1 0 13616 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_149
timestamp 1562078211
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_161
timestamp 1
transform 1 0 15824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_165
timestamp 1
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16376 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_169
timestamp 1562078211
transform 1 0 16560 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_181
timestamp 1562078211
transform 1 0 17664 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_193
timestamp 1562078211
transform 1 0 18768 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_205
timestamp 1562078211
transform 1 0 19872 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_217
timestamp 1
transform 1 0 20976 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1
transform 1 0 21344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_225
timestamp 1562078211
transform 1 0 21712 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_237
timestamp 1562078211
transform 1 0 22816 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_249
timestamp 1562078211
transform 1 0 23920 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_261
timestamp 1562078211
transform 1 0 25024 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_273
timestamp 1
transform 1 0 26128 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_277
timestamp 1
transform 1 0 26496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26680 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_281
timestamp 1562078211
transform 1 0 26864 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_293
timestamp 1562078211
transform 1 0 27968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_7_305
timestamp 1
transform 1 0 29072 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_313
timestamp 1
transform 1 0 29808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_324
timestamp 1
transform 1 0 30820 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_333
timestamp 1
transform 1 0 31648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1
transform 1 0 31832 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_343
timestamp 1562078211
transform 1 0 32568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_7_355
timestamp 1
transform 1 0 33672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_363
timestamp 1
transform 1 0 34408 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_367
timestamp 1
transform 1 0 34776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_369
timestamp 1
transform 1 0 34960 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_372
timestamp 1562078211
transform 1 0 35236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_7_384
timestamp 1
transform 1 0 36340 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_393
timestamp 1562078211
transform 1 0 37168 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_405
timestamp 1562078211
transform 1 0 38272 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_417
timestamp 1562078211
transform 1 0 39376 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_429
timestamp 1562078211
transform 1 0 40480 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_441
timestamp 1
transform 1 0 41584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_445
timestamp 1
transform 1 0 41952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1
transform 1 0 42136 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_449
timestamp 1562078211
transform 1 0 42320 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_461
timestamp 1562078211
transform 1 0 43424 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_473
timestamp 1
transform 1 0 44528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_523
timestamp 1562078211
transform 1 0 49128 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_535
timestamp 1
transform 1 0 50232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_537
timestamp 1
transform 1 0 50416 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_546
timestamp 1562078211
transform 1 0 51244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_558
timestamp 1
transform 1 0 52348 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_561
timestamp 1562078211
transform 1 0 52624 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_573
timestamp 1
transform 1 0 53728 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_577
timestamp 1
transform 1 0 54096 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_587
timestamp 1562078211
transform 1 0 55016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_599
timestamp 1562078211
transform 1 0 56120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_611
timestamp 1
transform 1 0 57224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1
transform 1 0 57592 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_617
timestamp 1562078211
transform 1 0 57776 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_629
timestamp 1
transform 1 0 58880 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_633
timestamp 1562078211
transform 1 0 59248 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_645
timestamp 1
transform 1 0 60352 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_649
timestamp 1562078211
transform 1 0 60720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_661
timestamp 1
transform 1 0 61824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_7_665
timestamp 1
transform 1 0 62192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_669
timestamp 1
transform 1 0 62560 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1
transform 1 0 62744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_7_673
timestamp 1
transform 1 0 62928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_677
timestamp 1
transform 1 0 63296 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_681
timestamp 1562078211
transform 1 0 63664 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_693
timestamp 1562078211
transform 1 0 64768 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_705
timestamp 1
transform 1 0 65872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_709
timestamp 1
transform 1 0 66240 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_713
timestamp 1562078211
transform 1 0 66608 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_725
timestamp 1
transform 1 0 67712 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1
transform 1 0 67896 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_729
timestamp 1562078211
transform 1 0 68080 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_743
timestamp 1562078211
transform 1 0 69368 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_755
timestamp 1562078211
transform 1 0 70472 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_767
timestamp 1562078211
transform 1 0 71576 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_779
timestamp 1
transform 1 0 72680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1
transform 1 0 73048 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_7_785
timestamp 1562078211
transform 1 0 73232 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_7_797
timestamp 1
transform 1 0 74336 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_3
timestamp 1562078211
transform 1 0 1288 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_15
timestamp 1562078211
transform 1 0 2392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_29
timestamp 1562078211
transform 1 0 3680 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_41
timestamp 1562078211
transform 1 0 4784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_57
timestamp 1562078211
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_69
timestamp 1562078211
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_85
timestamp 1562078211
transform 1 0 8832 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_97
timestamp 1562078211
transform 1 0 9936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1
transform 1 0 11040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp 1
transform 1 0 11224 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_113
timestamp 1562078211
transform 1 0 11408 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_125
timestamp 1562078211
transform 1 0 12512 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1
transform 1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13800 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_141
timestamp 1562078211
transform 1 0 13984 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_153
timestamp 1562078211
transform 1 0 15088 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1
transform 1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_167
timestamp 1
transform 1 0 16376 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_169
timestamp 1562078211
transform 1 0 16560 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_181
timestamp 1562078211
transform 1 0 17664 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_193
timestamp 1
transform 1 0 18768 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 18952 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_197
timestamp 1562078211
transform 1 0 19136 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_209
timestamp 1562078211
transform 1 0 20240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1
transform 1 0 21344 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_223
timestamp 1
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_225
timestamp 1562078211
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_237
timestamp 1562078211
transform 1 0 22816 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_249
timestamp 1
transform 1 0 23920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24104 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_253
timestamp 1562078211
transform 1 0 24288 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_265
timestamp 1562078211
transform 1 0 25392 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_277
timestamp 1
transform 1 0 26496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_279
timestamp 1
transform 1 0 26680 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_281
timestamp 1562078211
transform 1 0 26864 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_293
timestamp 1562078211
transform 1 0 27968 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_305
timestamp 1
transform 1 0 29072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1
transform 1 0 29256 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_309
timestamp 1562078211
transform 1 0 29440 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_321
timestamp 1562078211
transform 1 0 30544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_333
timestamp 1
transform 1 0 31648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_335
timestamp 1
transform 1 0 31832 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_337
timestamp 1562078211
transform 1 0 32016 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_349
timestamp 1562078211
transform 1 0 33120 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_361
timestamp 1
transform 1 0 34224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1
transform 1 0 34408 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_365
timestamp 1562078211
transform 1 0 34592 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_377
timestamp 1562078211
transform 1 0 35696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_389
timestamp 1
transform 1 0 36800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_391
timestamp 1
transform 1 0 36984 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_393
timestamp 1562078211
transform 1 0 37168 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_405
timestamp 1562078211
transform 1 0 38272 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_417
timestamp 1
transform 1 0 39376 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1
transform 1 0 39560 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_421
timestamp 1562078211
transform 1 0 39744 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_433
timestamp 1562078211
transform 1 0 40848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_445
timestamp 1
transform 1 0 41952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_447
timestamp 1
transform 1 0 42136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_449
timestamp 1
transform 1 0 42320 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_457
timestamp 1
transform 1 0 43056 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_465
timestamp 1
transform 1 0 43792 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_477
timestamp 1
transform 1 0 44896 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_479
timestamp 1
transform 1 0 45080 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_505
timestamp 1562078211
transform 1 0 47472 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_517
timestamp 1
transform 1 0 48576 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_529
timestamp 1
transform 1 0 49680 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1
transform 1 0 49864 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_557
timestamp 1
transform 1 0 52256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_559
timestamp 1
transform 1 0 52440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_585
timestamp 1
transform 1 0 54832 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1
transform 1 0 55016 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_613
timestamp 1
transform 1 0 57408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_615
timestamp 1
transform 1 0 57592 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_617
timestamp 1562078211
transform 1 0 57776 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_629
timestamp 1
transform 1 0 58880 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_8_639
timestamp 1
transform 1 0 59800 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1
transform 1 0 60168 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_645
timestamp 1
transform 1 0 60352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_8_655
timestamp 1
transform 1 0 61272 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_671
timestamp 1
transform 1 0 62744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_8_673
timestamp 1
transform 1 0 62928 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_677
timestamp 1
transform 1 0 63296 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_685
timestamp 1562078211
transform 1 0 64032 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_697
timestamp 1
transform 1 0 65136 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1
transform 1 0 65320 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_701
timestamp 1
transform 1 0 65504 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_709
timestamp 1
transform 1 0 66240 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_713
timestamp 1562078211
transform 1 0 66608 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_725
timestamp 1
transform 1 0 67712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_727
timestamp 1
transform 1 0 67896 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_729
timestamp 1562078211
transform 1 0 68080 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_743
timestamp 1562078211
transform 1 0 69368 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1
transform 1 0 70472 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_757
timestamp 1562078211
transform 1 0 70656 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_769
timestamp 1562078211
transform 1 0 71760 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_781
timestamp 1
transform 1 0 72864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_783
timestamp 1
transform 1 0 73048 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_8_785
timestamp 1562078211
transform 1 0 73232 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_8_797
timestamp 1
transform 1 0 74336 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_9_703
timestamp 1
transform 1 0 65688 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_713
timestamp 1562078211
transform 1 0 66608 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_725
timestamp 1562078211
transform 1 0 67712 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_9_737
timestamp 1
transform 1 0 68816 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_743
timestamp 1562078211
transform 1 0 69368 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_755
timestamp 1
transform 1 0 70472 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_757
timestamp 1562078211
transform 1 0 70656 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_769
timestamp 1562078211
transform 1 0 71760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_9_781
timestamp 1562078211
transform 1 0 72864 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_9_793
timestamp 1
transform 1 0 73968 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_703
timestamp 1
transform 1 0 65688 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_713
timestamp 1562078211
transform 1 0 66608 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_725
timestamp 1
transform 1 0 67712 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_727
timestamp 1
transform 1 0 67896 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_729
timestamp 1562078211
transform 1 0 68080 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_743
timestamp 1562078211
transform 1 0 69368 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_755
timestamp 1562078211
transform 1 0 70472 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_767
timestamp 1562078211
transform 1 0 71576 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_779
timestamp 1
transform 1 0 72680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_783
timestamp 1
transform 1 0 73048 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_10_785
timestamp 1562078211
transform 1 0 73232 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_10_797
timestamp 1
transform 1 0 74336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_705
timestamp 1
transform 1 0 65872 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_709
timestamp 1
transform 1 0 66240 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_713
timestamp 1562078211
transform 1 0 66608 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_725
timestamp 1562078211
transform 1 0 67712 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_11_737
timestamp 1
transform 1 0 68816 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_743
timestamp 1562078211
transform 1 0 69368 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_755
timestamp 1
transform 1 0 70472 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_757
timestamp 1562078211
transform 1 0 70656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_769
timestamp 1562078211
transform 1 0 71760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_11_781
timestamp 1562078211
transform 1 0 72864 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_11_793
timestamp 1
transform 1 0 73968 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_703
timestamp 1562078211
transform 1 0 65688 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_715
timestamp 1562078211
transform 1 0 66792 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_727
timestamp 1
transform 1 0 67896 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_729
timestamp 1562078211
transform 1 0 68080 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_741
timestamp 1562078211
transform 1 0 69184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_753
timestamp 1562078211
transform 1 0 70288 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_765
timestamp 1562078211
transform 1 0 71392 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_777
timestamp 1
transform 1 0 72496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_781
timestamp 1
transform 1 0 72864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_783
timestamp 1
transform 1 0 73048 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_12_785
timestamp 1562078211
transform 1 0 73232 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_12_797
timestamp 1
transform 1 0 74336 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_703
timestamp 1562078211
transform 1 0 65688 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_715
timestamp 1562078211
transform 1 0 66792 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_727
timestamp 1562078211
transform 1 0 67896 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_739
timestamp 1562078211
transform 1 0 69000 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_13_751
timestamp 1
transform 1 0 70104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_755
timestamp 1
transform 1 0 70472 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_757
timestamp 1562078211
transform 1 0 70656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_769
timestamp 1562078211
transform 1 0 71760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_13_781
timestamp 1562078211
transform 1 0 72864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_13_793
timestamp 1
transform 1 0 73968 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_703
timestamp 1562078211
transform 1 0 65688 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_715
timestamp 1562078211
transform 1 0 66792 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_727
timestamp 1
transform 1 0 67896 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_729
timestamp 1562078211
transform 1 0 68080 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_741
timestamp 1562078211
transform 1 0 69184 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_753
timestamp 1562078211
transform 1 0 70288 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_765
timestamp 1562078211
transform 1 0 71392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_777
timestamp 1
transform 1 0 72496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_781
timestamp 1
transform 1 0 72864 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_783
timestamp 1
transform 1 0 73048 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_14_785
timestamp 1562078211
transform 1 0 73232 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_14_797
timestamp 1
transform 1 0 74336 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_703
timestamp 1562078211
transform 1 0 65688 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_715
timestamp 1562078211
transform 1 0 66792 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_727
timestamp 1562078211
transform 1 0 67896 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_739
timestamp 1562078211
transform 1 0 69000 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_15_751
timestamp 1
transform 1 0 70104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_755
timestamp 1
transform 1 0 70472 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_757
timestamp 1562078211
transform 1 0 70656 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_769
timestamp 1562078211
transform 1 0 71760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_15_781
timestamp 1562078211
transform 1 0 72864 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_15_793
timestamp 1
transform 1 0 73968 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_703
timestamp 1562078211
transform 1 0 65688 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_715
timestamp 1562078211
transform 1 0 66792 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_727
timestamp 1
transform 1 0 67896 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_729
timestamp 1562078211
transform 1 0 68080 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_741
timestamp 1562078211
transform 1 0 69184 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_753
timestamp 1562078211
transform 1 0 70288 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_765
timestamp 1562078211
transform 1 0 71392 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_16_777
timestamp 1
transform 1 0 72496 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_781
timestamp 1
transform 1 0 72864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_783
timestamp 1
transform 1 0 73048 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_16_785
timestamp 1562078211
transform 1 0 73232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_16_797
timestamp 1
transform 1 0 74336 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_703
timestamp 1562078211
transform 1 0 65688 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_715
timestamp 1562078211
transform 1 0 66792 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_727
timestamp 1562078211
transform 1 0 67896 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_739
timestamp 1562078211
transform 1 0 69000 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_17_751
timestamp 1
transform 1 0 70104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_755
timestamp 1
transform 1 0 70472 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_757
timestamp 1562078211
transform 1 0 70656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_769
timestamp 1562078211
transform 1 0 71760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_17_781
timestamp 1562078211
transform 1 0 72864 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_17_793
timestamp 1
transform 1 0 73968 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_703
timestamp 1562078211
transform 1 0 65688 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_715
timestamp 1562078211
transform 1 0 66792 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_727
timestamp 1
transform 1 0 67896 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_729
timestamp 1562078211
transform 1 0 68080 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_741
timestamp 1562078211
transform 1 0 69184 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_753
timestamp 1562078211
transform 1 0 70288 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_765
timestamp 1562078211
transform 1 0 71392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_18_777
timestamp 1
transform 1 0 72496 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_781
timestamp 1
transform 1 0 72864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_783
timestamp 1
transform 1 0 73048 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_18_785
timestamp 1562078211
transform 1 0 73232 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_18_797
timestamp 1
transform 1 0 74336 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_703
timestamp 1562078211
transform 1 0 65688 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_715
timestamp 1562078211
transform 1 0 66792 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_727
timestamp 1562078211
transform 1 0 67896 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_739
timestamp 1562078211
transform 1 0 69000 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_19_751
timestamp 1
transform 1 0 70104 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_755
timestamp 1
transform 1 0 70472 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_757
timestamp 1562078211
transform 1 0 70656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_769
timestamp 1562078211
transform 1 0 71760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_19_781
timestamp 1562078211
transform 1 0 72864 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_19_793
timestamp 1
transform 1 0 73968 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_703
timestamp 1562078211
transform 1 0 65688 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_715
timestamp 1562078211
transform 1 0 66792 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_727
timestamp 1
transform 1 0 67896 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_729
timestamp 1562078211
transform 1 0 68080 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_741
timestamp 1562078211
transform 1 0 69184 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_753
timestamp 1562078211
transform 1 0 70288 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_765
timestamp 1562078211
transform 1 0 71392 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_20_777
timestamp 1
transform 1 0 72496 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_781
timestamp 1
transform 1 0 72864 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_783
timestamp 1
transform 1 0 73048 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_20_785
timestamp 1562078211
transform 1 0 73232 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_20_797
timestamp 1
transform 1 0 74336 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_703
timestamp 1562078211
transform 1 0 65688 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_715
timestamp 1562078211
transform 1 0 66792 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_727
timestamp 1562078211
transform 1 0 67896 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_739
timestamp 1562078211
transform 1 0 69000 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_21_751
timestamp 1
transform 1 0 70104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_755
timestamp 1
transform 1 0 70472 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_757
timestamp 1562078211
transform 1 0 70656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_769
timestamp 1562078211
transform 1 0 71760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_21_781
timestamp 1562078211
transform 1 0 72864 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_21_793
timestamp 1
transform 1 0 73968 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_703
timestamp 1562078211
transform 1 0 65688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_715
timestamp 1562078211
transform 1 0 66792 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_727
timestamp 1
transform 1 0 67896 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_729
timestamp 1562078211
transform 1 0 68080 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_741
timestamp 1562078211
transform 1 0 69184 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_753
timestamp 1562078211
transform 1 0 70288 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_765
timestamp 1562078211
transform 1 0 71392 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_22_777
timestamp 1
transform 1 0 72496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_781
timestamp 1
transform 1 0 72864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_783
timestamp 1
transform 1 0 73048 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_22_785
timestamp 1562078211
transform 1 0 73232 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_22_797
timestamp 1
transform 1 0 74336 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_703
timestamp 1562078211
transform 1 0 65688 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_715
timestamp 1562078211
transform 1 0 66792 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_727
timestamp 1562078211
transform 1 0 67896 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_739
timestamp 1562078211
transform 1 0 69000 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_23_751
timestamp 1
transform 1 0 70104 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_755
timestamp 1
transform 1 0 70472 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_757
timestamp 1562078211
transform 1 0 70656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_769
timestamp 1562078211
transform 1 0 71760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_23_781
timestamp 1562078211
transform 1 0 72864 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_23_793
timestamp 1
transform 1 0 73968 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_703
timestamp 1562078211
transform 1 0 65688 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_715
timestamp 1562078211
transform 1 0 66792 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_727
timestamp 1
transform 1 0 67896 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_729
timestamp 1562078211
transform 1 0 68080 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_741
timestamp 1562078211
transform 1 0 69184 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_753
timestamp 1562078211
transform 1 0 70288 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_765
timestamp 1562078211
transform 1 0 71392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_24_777
timestamp 1
transform 1 0 72496 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_781
timestamp 1
transform 1 0 72864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_783
timestamp 1
transform 1 0 73048 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_24_785
timestamp 1562078211
transform 1 0 73232 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_24_797
timestamp 1
transform 1 0 74336 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_703
timestamp 1562078211
transform 1 0 65688 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_715
timestamp 1562078211
transform 1 0 66792 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_727
timestamp 1562078211
transform 1 0 67896 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_739
timestamp 1562078211
transform 1 0 69000 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_25_751
timestamp 1
transform 1 0 70104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_755
timestamp 1
transform 1 0 70472 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_757
timestamp 1562078211
transform 1 0 70656 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_769
timestamp 1562078211
transform 1 0 71760 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_25_781
timestamp 1562078211
transform 1 0 72864 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_25_793
timestamp 1
transform 1 0 73968 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_703
timestamp 1562078211
transform 1 0 65688 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_715
timestamp 1562078211
transform 1 0 66792 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_727
timestamp 1
transform 1 0 67896 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_729
timestamp 1562078211
transform 1 0 68080 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_741
timestamp 1562078211
transform 1 0 69184 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_753
timestamp 1562078211
transform 1 0 70288 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_765
timestamp 1562078211
transform 1 0 71392 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_26_777
timestamp 1
transform 1 0 72496 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_781
timestamp 1
transform 1 0 72864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_783
timestamp 1
transform 1 0 73048 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_26_785
timestamp 1562078211
transform 1 0 73232 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_26_797
timestamp 1
transform 1 0 74336 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_703
timestamp 1562078211
transform 1 0 65688 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_715
timestamp 1562078211
transform 1 0 66792 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_727
timestamp 1562078211
transform 1 0 67896 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_739
timestamp 1562078211
transform 1 0 69000 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_27_751
timestamp 1
transform 1 0 70104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_755
timestamp 1
transform 1 0 70472 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_757
timestamp 1562078211
transform 1 0 70656 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_769
timestamp 1562078211
transform 1 0 71760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_27_781
timestamp 1562078211
transform 1 0 72864 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_27_793
timestamp 1
transform 1 0 73968 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_703
timestamp 1562078211
transform 1 0 65688 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_715
timestamp 1562078211
transform 1 0 66792 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_727
timestamp 1
transform 1 0 67896 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_729
timestamp 1562078211
transform 1 0 68080 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_741
timestamp 1562078211
transform 1 0 69184 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_753
timestamp 1562078211
transform 1 0 70288 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_765
timestamp 1562078211
transform 1 0 71392 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_28_777
timestamp 1
transform 1 0 72496 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_781
timestamp 1
transform 1 0 72864 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_783
timestamp 1
transform 1 0 73048 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_28_785
timestamp 1562078211
transform 1 0 73232 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_28_797
timestamp 1
transform 1 0 74336 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_703
timestamp 1562078211
transform 1 0 65688 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_715
timestamp 1562078211
transform 1 0 66792 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_727
timestamp 1562078211
transform 1 0 67896 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_739
timestamp 1562078211
transform 1 0 69000 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_29_751
timestamp 1
transform 1 0 70104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_755
timestamp 1
transform 1 0 70472 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_757
timestamp 1562078211
transform 1 0 70656 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_769
timestamp 1562078211
transform 1 0 71760 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_29_781
timestamp 1562078211
transform 1 0 72864 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_29_793
timestamp 1
transform 1 0 73968 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_703
timestamp 1562078211
transform 1 0 65688 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_715
timestamp 1562078211
transform 1 0 66792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_727
timestamp 1
transform 1 0 67896 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_729
timestamp 1562078211
transform 1 0 68080 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_741
timestamp 1562078211
transform 1 0 69184 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_753
timestamp 1562078211
transform 1 0 70288 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_765
timestamp 1562078211
transform 1 0 71392 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_30_777
timestamp 1
transform 1 0 72496 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_781
timestamp 1
transform 1 0 72864 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_783
timestamp 1
transform 1 0 73048 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_30_785
timestamp 1562078211
transform 1 0 73232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_30_797
timestamp 1
transform 1 0 74336 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_703
timestamp 1562078211
transform 1 0 65688 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_715
timestamp 1562078211
transform 1 0 66792 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_727
timestamp 1562078211
transform 1 0 67896 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_739
timestamp 1562078211
transform 1 0 69000 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_31_751
timestamp 1
transform 1 0 70104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_755
timestamp 1
transform 1 0 70472 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_757
timestamp 1562078211
transform 1 0 70656 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_769
timestamp 1562078211
transform 1 0 71760 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_31_781
timestamp 1562078211
transform 1 0 72864 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_31_793
timestamp 1
transform 1 0 73968 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_703
timestamp 1562078211
transform 1 0 65688 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_715
timestamp 1562078211
transform 1 0 66792 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_727
timestamp 1
transform 1 0 67896 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_729
timestamp 1562078211
transform 1 0 68080 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_741
timestamp 1562078211
transform 1 0 69184 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_753
timestamp 1562078211
transform 1 0 70288 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_765
timestamp 1562078211
transform 1 0 71392 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_32_777
timestamp 1
transform 1 0 72496 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_781
timestamp 1
transform 1 0 72864 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_783
timestamp 1
transform 1 0 73048 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_32_785
timestamp 1562078211
transform 1 0 73232 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_32_797
timestamp 1
transform 1 0 74336 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_703
timestamp 1562078211
transform 1 0 65688 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_715
timestamp 1562078211
transform 1 0 66792 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_727
timestamp 1562078211
transform 1 0 67896 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_739
timestamp 1562078211
transform 1 0 69000 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_33_751
timestamp 1
transform 1 0 70104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_755
timestamp 1
transform 1 0 70472 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_757
timestamp 1562078211
transform 1 0 70656 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_769
timestamp 1562078211
transform 1 0 71760 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_33_781
timestamp 1562078211
transform 1 0 72864 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_33_793
timestamp 1
transform 1 0 73968 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_703
timestamp 1562078211
transform 1 0 65688 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_715
timestamp 1562078211
transform 1 0 66792 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_727
timestamp 1
transform 1 0 67896 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_729
timestamp 1562078211
transform 1 0 68080 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_741
timestamp 1562078211
transform 1 0 69184 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_753
timestamp 1562078211
transform 1 0 70288 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_765
timestamp 1562078211
transform 1 0 71392 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_777
timestamp 1
transform 1 0 72496 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_781
timestamp 1
transform 1 0 72864 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_783
timestamp 1
transform 1 0 73048 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_34_785
timestamp 1562078211
transform 1 0 73232 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_34_797
timestamp 1
transform 1 0 74336 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_703
timestamp 1562078211
transform 1 0 65688 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_715
timestamp 1562078211
transform 1 0 66792 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_727
timestamp 1562078211
transform 1 0 67896 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_739
timestamp 1562078211
transform 1 0 69000 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_35_751
timestamp 1
transform 1 0 70104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_755
timestamp 1
transform 1 0 70472 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_757
timestamp 1562078211
transform 1 0 70656 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_769
timestamp 1562078211
transform 1 0 71760 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_35_781
timestamp 1562078211
transform 1 0 72864 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_35_793
timestamp 1
transform 1 0 73968 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_703
timestamp 1562078211
transform 1 0 65688 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_715
timestamp 1562078211
transform 1 0 66792 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_727
timestamp 1
transform 1 0 67896 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_729
timestamp 1562078211
transform 1 0 68080 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_741
timestamp 1562078211
transform 1 0 69184 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_753
timestamp 1562078211
transform 1 0 70288 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_765
timestamp 1562078211
transform 1 0 71392 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_36_777
timestamp 1
transform 1 0 72496 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_781
timestamp 1
transform 1 0 72864 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_783
timestamp 1
transform 1 0 73048 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_36_785
timestamp 1562078211
transform 1 0 73232 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_36_797
timestamp 1
transform 1 0 74336 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_703
timestamp 1562078211
transform 1 0 65688 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_715
timestamp 1562078211
transform 1 0 66792 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_727
timestamp 1562078211
transform 1 0 67896 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_739
timestamp 1562078211
transform 1 0 69000 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_37_751
timestamp 1
transform 1 0 70104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_755
timestamp 1
transform 1 0 70472 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_757
timestamp 1562078211
transform 1 0 70656 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_769
timestamp 1562078211
transform 1 0 71760 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_37_781
timestamp 1562078211
transform 1 0 72864 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_37_793
timestamp 1
transform 1 0 73968 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_703
timestamp 1562078211
transform 1 0 65688 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_715
timestamp 1562078211
transform 1 0 66792 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_727
timestamp 1
transform 1 0 67896 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_729
timestamp 1562078211
transform 1 0 68080 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_741
timestamp 1562078211
transform 1 0 69184 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_753
timestamp 1562078211
transform 1 0 70288 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_765
timestamp 1562078211
transform 1 0 71392 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_38_777
timestamp 1
transform 1 0 72496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_781
timestamp 1
transform 1 0 72864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_783
timestamp 1
transform 1 0 73048 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_38_785
timestamp 1562078211
transform 1 0 73232 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_38_797
timestamp 1
transform 1 0 74336 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_711
timestamp 1562078211
transform 1 0 66424 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_723
timestamp 1562078211
transform 1 0 67528 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_735
timestamp 1562078211
transform 1 0 68632 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_39_747
timestamp 1
transform 1 0 69736 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_755
timestamp 1
transform 1 0 70472 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_757
timestamp 1562078211
transform 1 0 70656 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_769
timestamp 1562078211
transform 1 0 71760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_39_781
timestamp 1562078211
transform 1 0 72864 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_39_793
timestamp 1
transform 1 0 73968 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_721
timestamp 1
transform 1 0 67344 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_725
timestamp 1
transform 1 0 67712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_727
timestamp 1
transform 1 0 67896 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_729
timestamp 1562078211
transform 1 0 68080 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_741
timestamp 1562078211
transform 1 0 69184 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_753
timestamp 1562078211
transform 1 0 70288 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_765
timestamp 1562078211
transform 1 0 71392 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_40_777
timestamp 1
transform 1 0 72496 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_781
timestamp 1
transform 1 0 72864 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_783
timestamp 1
transform 1 0 73048 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_40_785
timestamp 1562078211
transform 1 0 73232 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_40_797
timestamp 1
transform 1 0 74336 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_727
timestamp 1562078211
transform 1 0 67896 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_739
timestamp 1562078211
transform 1 0 69000 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_41_751
timestamp 1
transform 1 0 70104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_755
timestamp 1
transform 1 0 70472 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_757
timestamp 1562078211
transform 1 0 70656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_769
timestamp 1562078211
transform 1 0 71760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_41_781
timestamp 1562078211
transform 1 0 72864 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_41_793
timestamp 1
transform 1 0 73968 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_721
timestamp 1
transform 1 0 67344 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_725
timestamp 1
transform 1 0 67712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_727
timestamp 1
transform 1 0 67896 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_729
timestamp 1562078211
transform 1 0 68080 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_741
timestamp 1562078211
transform 1 0 69184 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_753
timestamp 1562078211
transform 1 0 70288 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_765
timestamp 1562078211
transform 1 0 71392 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_777
timestamp 1
transform 1 0 72496 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_781
timestamp 1
transform 1 0 72864 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_783
timestamp 1
transform 1 0 73048 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_42_785
timestamp 1562078211
transform 1 0 73232 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_42_797
timestamp 1
transform 1 0 74336 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_715
timestamp 1562078211
transform 1 0 66792 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_727
timestamp 1562078211
transform 1 0 67896 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_739
timestamp 1562078211
transform 1 0 69000 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_43_751
timestamp 1
transform 1 0 70104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_755
timestamp 1
transform 1 0 70472 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_757
timestamp 1562078211
transform 1 0 70656 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_769
timestamp 1562078211
transform 1 0 71760 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_43_781
timestamp 1562078211
transform 1 0 72864 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_43_793
timestamp 1
transform 1 0 73968 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_711
timestamp 1562078211
transform 1 0 66424 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_44_723
timestamp 1
transform 1 0 67528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_727
timestamp 1
transform 1 0 67896 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_729
timestamp 1562078211
transform 1 0 68080 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_741
timestamp 1562078211
transform 1 0 69184 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_753
timestamp 1562078211
transform 1 0 70288 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_765
timestamp 1562078211
transform 1 0 71392 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_44_777
timestamp 1
transform 1 0 72496 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_781
timestamp 1
transform 1 0 72864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_783
timestamp 1
transform 1 0 73048 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_44_785
timestamp 1562078211
transform 1 0 73232 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_44_797
timestamp 1
transform 1 0 74336 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_703
timestamp 1562078211
transform 1 0 65688 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_715
timestamp 1562078211
transform 1 0 66792 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_727
timestamp 1562078211
transform 1 0 67896 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_739
timestamp 1562078211
transform 1 0 69000 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_45_751
timestamp 1
transform 1 0 70104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_755
timestamp 1
transform 1 0 70472 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_757
timestamp 1562078211
transform 1 0 70656 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_769
timestamp 1562078211
transform 1 0 71760 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_45_781
timestamp 1562078211
transform 1 0 72864 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_45_793
timestamp 1
transform 1 0 73968 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_711
timestamp 1562078211
transform 1 0 66424 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_46_723
timestamp 1
transform 1 0 67528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_727
timestamp 1
transform 1 0 67896 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_729
timestamp 1562078211
transform 1 0 68080 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_741
timestamp 1562078211
transform 1 0 69184 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_753
timestamp 1562078211
transform 1 0 70288 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_765
timestamp 1562078211
transform 1 0 71392 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_46_777
timestamp 1
transform 1 0 72496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_781
timestamp 1
transform 1 0 72864 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_783
timestamp 1
transform 1 0 73048 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_46_785
timestamp 1562078211
transform 1 0 73232 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_46_797
timestamp 1
transform 1 0 74336 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_719
timestamp 1562078211
transform 1 0 67160 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_731
timestamp 1562078211
transform 1 0 68264 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_743
timestamp 1562078211
transform 1 0 69368 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_755
timestamp 1
transform 1 0 70472 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_757
timestamp 1562078211
transform 1 0 70656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_769
timestamp 1562078211
transform 1 0 71760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_47_781
timestamp 1562078211
transform 1 0 72864 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_47_793
timestamp 1
transform 1 0 73968 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_711
timestamp 1562078211
transform 1 0 66424 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_48_723
timestamp 1
transform 1 0 67528 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_727
timestamp 1
transform 1 0 67896 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_729
timestamp 1562078211
transform 1 0 68080 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_741
timestamp 1562078211
transform 1 0 69184 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_753
timestamp 1562078211
transform 1 0 70288 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_765
timestamp 1562078211
transform 1 0 71392 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_48_777
timestamp 1
transform 1 0 72496 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_781
timestamp 1
transform 1 0 72864 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_783
timestamp 1
transform 1 0 73048 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_48_785
timestamp 1562078211
transform 1 0 73232 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_48_797
timestamp 1
transform 1 0 74336 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_711
timestamp 1562078211
transform 1 0 66424 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_723
timestamp 1562078211
transform 1 0 67528 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_735
timestamp 1562078211
transform 1 0 68632 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_49_747
timestamp 1
transform 1 0 69736 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_755
timestamp 1
transform 1 0 70472 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_757
timestamp 1562078211
transform 1 0 70656 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_769
timestamp 1562078211
transform 1 0 71760 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_49_781
timestamp 1562078211
transform 1 0 72864 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_49_793
timestamp 1
transform 1 0 73968 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_723
timestamp 1
transform 1 0 67528 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_727
timestamp 1
transform 1 0 67896 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_729
timestamp 1562078211
transform 1 0 68080 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_741
timestamp 1562078211
transform 1 0 69184 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_753
timestamp 1562078211
transform 1 0 70288 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_765
timestamp 1562078211
transform 1 0 71392 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_50_777
timestamp 1
transform 1 0 72496 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_781
timestamp 1
transform 1 0 72864 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_783
timestamp 1
transform 1 0 73048 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_50_785
timestamp 1562078211
transform 1 0 73232 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_50_797
timestamp 1
transform 1 0 74336 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_703
timestamp 1562078211
transform 1 0 65688 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_715
timestamp 1562078211
transform 1 0 66792 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_727
timestamp 1562078211
transform 1 0 67896 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_739
timestamp 1562078211
transform 1 0 69000 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_51_751
timestamp 1
transform 1 0 70104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_755
timestamp 1
transform 1 0 70472 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_757
timestamp 1562078211
transform 1 0 70656 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_769
timestamp 1562078211
transform 1 0 71760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_51_781
timestamp 1562078211
transform 1 0 72864 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_51_793
timestamp 1
transform 1 0 73968 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_711
timestamp 1562078211
transform 1 0 66424 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_723
timestamp 1
transform 1 0 67528 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_727
timestamp 1
transform 1 0 67896 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_729
timestamp 1562078211
transform 1 0 68080 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_741
timestamp 1562078211
transform 1 0 69184 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_753
timestamp 1562078211
transform 1 0 70288 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_765
timestamp 1562078211
transform 1 0 71392 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_777
timestamp 1
transform 1 0 72496 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_781
timestamp 1
transform 1 0 72864 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_783
timestamp 1
transform 1 0 73048 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_52_785
timestamp 1562078211
transform 1 0 73232 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_52_797
timestamp 1
transform 1 0 74336 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_703
timestamp 1562078211
transform 1 0 65688 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_715
timestamp 1562078211
transform 1 0 66792 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_727
timestamp 1562078211
transform 1 0 67896 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_739
timestamp 1562078211
transform 1 0 69000 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_53_751
timestamp 1
transform 1 0 70104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_755
timestamp 1
transform 1 0 70472 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_757
timestamp 1562078211
transform 1 0 70656 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_769
timestamp 1562078211
transform 1 0 71760 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_53_781
timestamp 1562078211
transform 1 0 72864 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_53_793
timestamp 1
transform 1 0 73968 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_711
timestamp 1562078211
transform 1 0 66424 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_723
timestamp 1
transform 1 0 67528 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_727
timestamp 1
transform 1 0 67896 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_729
timestamp 1562078211
transform 1 0 68080 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_741
timestamp 1562078211
transform 1 0 69184 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_753
timestamp 1562078211
transform 1 0 70288 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_765
timestamp 1562078211
transform 1 0 71392 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_777
timestamp 1
transform 1 0 72496 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_781
timestamp 1
transform 1 0 72864 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_783
timestamp 1
transform 1 0 73048 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_54_785
timestamp 1562078211
transform 1 0 73232 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_54_797
timestamp 1
transform 1 0 74336 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_703
timestamp 1562078211
transform 1 0 65688 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_715
timestamp 1562078211
transform 1 0 66792 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_727
timestamp 1562078211
transform 1 0 67896 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_739
timestamp 1562078211
transform 1 0 69000 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_55_751
timestamp 1
transform 1 0 70104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_755
timestamp 1
transform 1 0 70472 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_757
timestamp 1562078211
transform 1 0 70656 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_769
timestamp 1562078211
transform 1 0 71760 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_55_781
timestamp 1562078211
transform 1 0 72864 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_55_793
timestamp 1
transform 1 0 73968 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_711
timestamp 1562078211
transform 1 0 66424 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_56_723
timestamp 1
transform 1 0 67528 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_727
timestamp 1
transform 1 0 67896 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_729
timestamp 1562078211
transform 1 0 68080 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_741
timestamp 1562078211
transform 1 0 69184 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_753
timestamp 1562078211
transform 1 0 70288 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_765
timestamp 1562078211
transform 1 0 71392 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_56_777
timestamp 1
transform 1 0 72496 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_781
timestamp 1
transform 1 0 72864 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_783
timestamp 1
transform 1 0 73048 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_56_785
timestamp 1562078211
transform 1 0 73232 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_56_797
timestamp 1
transform 1 0 74336 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_703
timestamp 1562078211
transform 1 0 65688 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_715
timestamp 1562078211
transform 1 0 66792 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_727
timestamp 1562078211
transform 1 0 67896 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_739
timestamp 1562078211
transform 1 0 69000 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_57_751
timestamp 1
transform 1 0 70104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_755
timestamp 1
transform 1 0 70472 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_757
timestamp 1562078211
transform 1 0 70656 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_769
timestamp 1562078211
transform 1 0 71760 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_57_781
timestamp 1562078211
transform 1 0 72864 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_57_793
timestamp 1
transform 1 0 73968 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_711
timestamp 1562078211
transform 1 0 66424 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_723
timestamp 1
transform 1 0 67528 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_727
timestamp 1
transform 1 0 67896 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_729
timestamp 1562078211
transform 1 0 68080 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_741
timestamp 1562078211
transform 1 0 69184 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_753
timestamp 1562078211
transform 1 0 70288 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_765
timestamp 1562078211
transform 1 0 71392 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_777
timestamp 1
transform 1 0 72496 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_781
timestamp 1
transform 1 0 72864 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_783
timestamp 1
transform 1 0 73048 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_58_785
timestamp 1562078211
transform 1 0 73232 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_58_797
timestamp 1
transform 1 0 74336 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_703
timestamp 1562078211
transform 1 0 65688 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_715
timestamp 1562078211
transform 1 0 66792 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_727
timestamp 1562078211
transform 1 0 67896 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_739
timestamp 1562078211
transform 1 0 69000 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_59_751
timestamp 1
transform 1 0 70104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_755
timestamp 1
transform 1 0 70472 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_757
timestamp 1562078211
transform 1 0 70656 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_769
timestamp 1562078211
transform 1 0 71760 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_59_781
timestamp 1562078211
transform 1 0 72864 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_59_793
timestamp 1
transform 1 0 73968 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_711
timestamp 1562078211
transform 1 0 66424 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_723
timestamp 1
transform 1 0 67528 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_727
timestamp 1
transform 1 0 67896 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_729
timestamp 1562078211
transform 1 0 68080 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_741
timestamp 1562078211
transform 1 0 69184 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_753
timestamp 1562078211
transform 1 0 70288 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_765
timestamp 1562078211
transform 1 0 71392 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_777
timestamp 1
transform 1 0 72496 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_781
timestamp 1
transform 1 0 72864 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_783
timestamp 1
transform 1 0 73048 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_60_785
timestamp 1562078211
transform 1 0 73232 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_60_797
timestamp 1
transform 1 0 74336 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_711
timestamp 1562078211
transform 1 0 66424 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_723
timestamp 1562078211
transform 1 0 67528 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_735
timestamp 1562078211
transform 1 0 68632 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_61_747
timestamp 1
transform 1 0 69736 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_755
timestamp 1
transform 1 0 70472 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_757
timestamp 1562078211
transform 1 0 70656 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_769
timestamp 1562078211
transform 1 0 71760 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_61_781
timestamp 1562078211
transform 1 0 72864 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_61_793
timestamp 1
transform 1 0 73968 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_719
timestamp 1
transform 1 0 67160 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_727
timestamp 1
transform 1 0 67896 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_729
timestamp 1562078211
transform 1 0 68080 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_741
timestamp 1562078211
transform 1 0 69184 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_753
timestamp 1562078211
transform 1 0 70288 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_765
timestamp 1562078211
transform 1 0 71392 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_62_777
timestamp 1
transform 1 0 72496 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_781
timestamp 1
transform 1 0 72864 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_783
timestamp 1
transform 1 0 73048 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_62_785
timestamp 1562078211
transform 1 0 73232 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_62_797
timestamp 1
transform 1 0 74336 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_723
timestamp 1562078211
transform 1 0 67528 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_735
timestamp 1562078211
transform 1 0 68632 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_63_747
timestamp 1
transform 1 0 69736 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_755
timestamp 1
transform 1 0 70472 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_757
timestamp 1562078211
transform 1 0 70656 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_769
timestamp 1562078211
transform 1 0 71760 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_63_781
timestamp 1562078211
transform 1 0 72864 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_63_793
timestamp 1
transform 1 0 73968 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_711
timestamp 1562078211
transform 1 0 66424 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_64_723
timestamp 1
transform 1 0 67528 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_727
timestamp 1
transform 1 0 67896 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_729
timestamp 1562078211
transform 1 0 68080 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_741
timestamp 1562078211
transform 1 0 69184 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_753
timestamp 1562078211
transform 1 0 70288 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_765
timestamp 1562078211
transform 1 0 71392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_64_777
timestamp 1
transform 1 0 72496 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_781
timestamp 1
transform 1 0 72864 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_783
timestamp 1
transform 1 0 73048 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_64_785
timestamp 1562078211
transform 1 0 73232 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_64_797
timestamp 1
transform 1 0 74336 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_703
timestamp 1562078211
transform 1 0 65688 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_715
timestamp 1562078211
transform 1 0 66792 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_727
timestamp 1562078211
transform 1 0 67896 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_739
timestamp 1562078211
transform 1 0 69000 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_65_751
timestamp 1
transform 1 0 70104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_755
timestamp 1
transform 1 0 70472 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_757
timestamp 1562078211
transform 1 0 70656 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_769
timestamp 1562078211
transform 1 0 71760 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_65_781
timestamp 1562078211
transform 1 0 72864 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_65_793
timestamp 1
transform 1 0 73968 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_703
timestamp 1562078211
transform 1 0 65688 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_715
timestamp 1562078211
transform 1 0 66792 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_727
timestamp 1
transform 1 0 67896 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_729
timestamp 1562078211
transform 1 0 68080 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_741
timestamp 1562078211
transform 1 0 69184 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_753
timestamp 1562078211
transform 1 0 70288 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_765
timestamp 1562078211
transform 1 0 71392 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_66_777
timestamp 1
transform 1 0 72496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_781
timestamp 1
transform 1 0 72864 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_783
timestamp 1
transform 1 0 73048 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_66_785
timestamp 1562078211
transform 1 0 73232 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_66_797
timestamp 1
transform 1 0 74336 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_711
timestamp 1562078211
transform 1 0 66424 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_723
timestamp 1562078211
transform 1 0 67528 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_735
timestamp 1562078211
transform 1 0 68632 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_67_747
timestamp 1
transform 1 0 69736 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_755
timestamp 1
transform 1 0 70472 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_757
timestamp 1562078211
transform 1 0 70656 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_769
timestamp 1562078211
transform 1 0 71760 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_67_781
timestamp 1562078211
transform 1 0 72864 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_67_793
timestamp 1
transform 1 0 73968 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_711
timestamp 1562078211
transform 1 0 66424 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_68_723
timestamp 1
transform 1 0 67528 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_727
timestamp 1
transform 1 0 67896 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_729
timestamp 1562078211
transform 1 0 68080 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_741
timestamp 1562078211
transform 1 0 69184 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_753
timestamp 1562078211
transform 1 0 70288 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_765
timestamp 1562078211
transform 1 0 71392 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_68_777
timestamp 1
transform 1 0 72496 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_781
timestamp 1
transform 1 0 72864 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_783
timestamp 1
transform 1 0 73048 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_68_785
timestamp 1562078211
transform 1 0 73232 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_68_797
timestamp 1
transform 1 0 74336 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_703
timestamp 1562078211
transform 1 0 65688 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_715
timestamp 1562078211
transform 1 0 66792 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_727
timestamp 1562078211
transform 1 0 67896 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_739
timestamp 1562078211
transform 1 0 69000 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_69_751
timestamp 1
transform 1 0 70104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_755
timestamp 1
transform 1 0 70472 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_757
timestamp 1562078211
transform 1 0 70656 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_769
timestamp 1562078211
transform 1 0 71760 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_69_781
timestamp 1562078211
transform 1 0 72864 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_69_793
timestamp 1
transform 1 0 73968 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_711
timestamp 1562078211
transform 1 0 66424 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_723
timestamp 1
transform 1 0 67528 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_727
timestamp 1
transform 1 0 67896 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_729
timestamp 1562078211
transform 1 0 68080 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_741
timestamp 1562078211
transform 1 0 69184 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_753
timestamp 1562078211
transform 1 0 70288 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_765
timestamp 1562078211
transform 1 0 71392 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_777
timestamp 1
transform 1 0 72496 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_781
timestamp 1
transform 1 0 72864 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_783
timestamp 1
transform 1 0 73048 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_70_785
timestamp 1562078211
transform 1 0 73232 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_70_797
timestamp 1
transform 1 0 74336 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_703
timestamp 1562078211
transform 1 0 65688 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_715
timestamp 1562078211
transform 1 0 66792 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_727
timestamp 1562078211
transform 1 0 67896 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_739
timestamp 1562078211
transform 1 0 69000 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_71_751
timestamp 1
transform 1 0 70104 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_755
timestamp 1
transform 1 0 70472 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_757
timestamp 1562078211
transform 1 0 70656 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_769
timestamp 1562078211
transform 1 0 71760 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_71_781
timestamp 1562078211
transform 1 0 72864 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_71_793
timestamp 1
transform 1 0 73968 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_703
timestamp 1
transform 1 0 65688 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_719
timestamp 1
transform 1 0 67160 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_727
timestamp 1
transform 1 0 67896 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_729
timestamp 1562078211
transform 1 0 68080 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_741
timestamp 1562078211
transform 1 0 69184 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_753
timestamp 1562078211
transform 1 0 70288 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_765
timestamp 1562078211
transform 1 0 71392 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_777
timestamp 1
transform 1 0 72496 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_781
timestamp 1
transform 1 0 72864 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_783
timestamp 1
transform 1 0 73048 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_72_785
timestamp 1562078211
transform 1 0 73232 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_72_797
timestamp 1
transform 1 0 74336 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_703
timestamp 1562078211
transform 1 0 65688 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_715
timestamp 1562078211
transform 1 0 66792 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_727
timestamp 1562078211
transform 1 0 67896 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_739
timestamp 1562078211
transform 1 0 69000 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_73_751
timestamp 1
transform 1 0 70104 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_755
timestamp 1
transform 1 0 70472 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_757
timestamp 1562078211
transform 1 0 70656 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_769
timestamp 1562078211
transform 1 0 71760 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_73_781
timestamp 1562078211
transform 1 0 72864 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_73_793
timestamp 1
transform 1 0 73968 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_703
timestamp 1
transform 1 0 65688 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_711
timestamp 1
transform 1 0 66424 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_713
timestamp 1
transform 1 0 66608 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_722
timestamp 1
transform 1 0 67436 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_726
timestamp 1
transform 1 0 67804 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_729
timestamp 1562078211
transform 1 0 68080 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_741
timestamp 1562078211
transform 1 0 69184 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_753
timestamp 1562078211
transform 1 0 70288 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_765
timestamp 1562078211
transform 1 0 71392 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_74_777
timestamp 1
transform 1 0 72496 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_781
timestamp 1
transform 1 0 72864 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_783
timestamp 1
transform 1 0 73048 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_74_785
timestamp 1562078211
transform 1 0 73232 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_74_797
timestamp 1
transform 1 0 74336 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_703
timestamp 1562078211
transform 1 0 65688 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_715
timestamp 1562078211
transform 1 0 66792 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_727
timestamp 1562078211
transform 1 0 67896 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_739
timestamp 1562078211
transform 1 0 69000 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_751
timestamp 1
transform 1 0 70104 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_755
timestamp 1
transform 1 0 70472 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_757
timestamp 1562078211
transform 1 0 70656 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_769
timestamp 1562078211
transform 1 0 71760 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_75_781
timestamp 1562078211
transform 1 0 72864 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_75_793
timestamp 1
transform 1 0 73968 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_706
timestamp 1562078211
transform 1 0 65964 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_76_718
timestamp 1
transform 1 0 67068 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_726
timestamp 1
transform 1 0 67804 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_737
timestamp 1562078211
transform 1 0 68816 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_749
timestamp 1562078211
transform 1 0 69920 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_761
timestamp 1562078211
transform 1 0 71024 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_76_773
timestamp 1
transform 1 0 72128 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_781
timestamp 1
transform 1 0 72864 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_783
timestamp 1
transform 1 0 73048 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_76_785
timestamp 1562078211
transform 1 0 73232 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_76_797
timestamp 1
transform 1 0 74336 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_703
timestamp 1562078211
transform 1 0 65688 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_715
timestamp 1562078211
transform 1 0 66792 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_727
timestamp 1562078211
transform 1 0 67896 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_739
timestamp 1562078211
transform 1 0 69000 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_77_751
timestamp 1
transform 1 0 70104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_755
timestamp 1
transform 1 0 70472 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_757
timestamp 1562078211
transform 1 0 70656 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_769
timestamp 1562078211
transform 1 0 71760 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_77_781
timestamp 1562078211
transform 1 0 72864 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_77_793
timestamp 1
transform 1 0 73968 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_706
timestamp 1562078211
transform 1 0 65964 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_78_718
timestamp 1
transform 1 0 67068 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_726
timestamp 1
transform 1 0 67804 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_729
timestamp 1562078211
transform 1 0 68080 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_741
timestamp 1562078211
transform 1 0 69184 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_753
timestamp 1562078211
transform 1 0 70288 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_765
timestamp 1562078211
transform 1 0 71392 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_78_777
timestamp 1
transform 1 0 72496 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_781
timestamp 1
transform 1 0 72864 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_783
timestamp 1
transform 1 0 73048 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_78_785
timestamp 1562078211
transform 1 0 73232 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_78_797
timestamp 1
transform 1 0 74336 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_703
timestamp 1562078211
transform 1 0 65688 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_715
timestamp 1562078211
transform 1 0 66792 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_727
timestamp 1562078211
transform 1 0 67896 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_739
timestamp 1562078211
transform 1 0 69000 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_79_751
timestamp 1
transform 1 0 70104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_755
timestamp 1
transform 1 0 70472 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_757
timestamp 1562078211
transform 1 0 70656 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_769
timestamp 1562078211
transform 1 0 71760 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_79_781
timestamp 1562078211
transform 1 0 72864 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_79_793
timestamp 1
transform 1 0 73968 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_703
timestamp 1562078211
transform 1 0 65688 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_715
timestamp 1562078211
transform 1 0 66792 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_727
timestamp 1
transform 1 0 67896 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_729
timestamp 1562078211
transform 1 0 68080 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_741
timestamp 1562078211
transform 1 0 69184 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_753
timestamp 1562078211
transform 1 0 70288 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_765
timestamp 1562078211
transform 1 0 71392 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_777
timestamp 1
transform 1 0 72496 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_781
timestamp 1
transform 1 0 72864 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_783
timestamp 1
transform 1 0 73048 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_80_785
timestamp 1562078211
transform 1 0 73232 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_80_797
timestamp 1
transform 1 0 74336 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_703
timestamp 1562078211
transform 1 0 65688 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_715
timestamp 1562078211
transform 1 0 66792 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_727
timestamp 1562078211
transform 1 0 67896 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_739
timestamp 1562078211
transform 1 0 69000 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_81_751
timestamp 1
transform 1 0 70104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_755
timestamp 1
transform 1 0 70472 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_757
timestamp 1562078211
transform 1 0 70656 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_769
timestamp 1562078211
transform 1 0 71760 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_81_781
timestamp 1562078211
transform 1 0 72864 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_81_793
timestamp 1
transform 1 0 73968 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_703
timestamp 1562078211
transform 1 0 65688 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_715
timestamp 1562078211
transform 1 0 66792 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_727
timestamp 1
transform 1 0 67896 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_729
timestamp 1562078211
transform 1 0 68080 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_741
timestamp 1562078211
transform 1 0 69184 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_753
timestamp 1562078211
transform 1 0 70288 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_765
timestamp 1562078211
transform 1 0 71392 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_82_777
timestamp 1
transform 1 0 72496 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_781
timestamp 1
transform 1 0 72864 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_783
timestamp 1
transform 1 0 73048 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_82_785
timestamp 1562078211
transform 1 0 73232 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_82_797
timestamp 1
transform 1 0 74336 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_83_703
timestamp 1562078211
transform 1 0 65688 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_83_715
timestamp 1562078211
transform 1 0 66792 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_83_727
timestamp 1562078211
transform 1 0 67896 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_83_739
timestamp 1562078211
transform 1 0 69000 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_83_751
timestamp 1
transform 1 0 70104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_755
timestamp 1
transform 1 0 70472 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_83_757
timestamp 1562078211
transform 1 0 70656 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_83_769
timestamp 1562078211
transform 1 0 71760 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_83_781
timestamp 1562078211
transform 1 0 72864 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_83_793
timestamp 1
transform 1 0 73968 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_84_709
timestamp 1562078211
transform 1 0 66240 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_84_721
timestamp 1
transform 1 0 67344 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_725
timestamp 1
transform 1 0 67712 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_727
timestamp 1
transform 1 0 67896 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_84_729
timestamp 1562078211
transform 1 0 68080 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_84_741
timestamp 1562078211
transform 1 0 69184 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_84_753
timestamp 1562078211
transform 1 0 70288 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_84_765
timestamp 1562078211
transform 1 0 71392 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_84_777
timestamp 1
transform 1 0 72496 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_781
timestamp 1
transform 1 0 72864 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_783
timestamp 1
transform 1 0 73048 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_84_785
timestamp 1562078211
transform 1 0 73232 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_84_797
timestamp 1
transform 1 0 74336 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_85_703
timestamp 1562078211
transform 1 0 65688 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_85_715
timestamp 1562078211
transform 1 0 66792 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_85_727
timestamp 1562078211
transform 1 0 67896 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_85_739
timestamp 1562078211
transform 1 0 69000 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_85_751
timestamp 1
transform 1 0 70104 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_755
timestamp 1
transform 1 0 70472 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_85_757
timestamp 1562078211
transform 1 0 70656 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_85_769
timestamp 1562078211
transform 1 0 71760 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_85_781
timestamp 1562078211
transform 1 0 72864 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_85_793
timestamp 1
transform 1 0 73968 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_86_703
timestamp 1562078211
transform 1 0 65688 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_86_715
timestamp 1562078211
transform 1 0 66792 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_727
timestamp 1
transform 1 0 67896 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_86_729
timestamp 1562078211
transform 1 0 68080 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_86_741
timestamp 1562078211
transform 1 0 69184 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_86_753
timestamp 1562078211
transform 1 0 70288 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_86_765
timestamp 1562078211
transform 1 0 71392 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_86_777
timestamp 1
transform 1 0 72496 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_781
timestamp 1
transform 1 0 72864 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_783
timestamp 1
transform 1 0 73048 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_86_785
timestamp 1562078211
transform 1 0 73232 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_86_797
timestamp 1
transform 1 0 74336 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_87_703
timestamp 1562078211
transform 1 0 65688 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_87_715
timestamp 1562078211
transform 1 0 66792 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_87_727
timestamp 1562078211
transform 1 0 67896 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_87_739
timestamp 1562078211
transform 1 0 69000 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_87_751
timestamp 1
transform 1 0 70104 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_755
timestamp 1
transform 1 0 70472 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_87_757
timestamp 1562078211
transform 1 0 70656 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_87_769
timestamp 1562078211
transform 1 0 71760 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_87_781
timestamp 1562078211
transform 1 0 72864 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_87_793
timestamp 1
transform 1 0 73968 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_88_706
timestamp 1562078211
transform 1 0 65964 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_88_718
timestamp 1
transform 1 0 67068 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_726
timestamp 1
transform 1 0 67804 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_88_729
timestamp 1562078211
transform 1 0 68080 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_88_741
timestamp 1562078211
transform 1 0 69184 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_88_753
timestamp 1562078211
transform 1 0 70288 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_88_765
timestamp 1562078211
transform 1 0 71392 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_88_777
timestamp 1
transform 1 0 72496 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_781
timestamp 1
transform 1 0 72864 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_783
timestamp 1
transform 1 0 73048 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_88_785
timestamp 1562078211
transform 1 0 73232 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_88_797
timestamp 1
transform 1 0 74336 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_89_706
timestamp 1562078211
transform 1 0 65964 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_89_718
timestamp 1562078211
transform 1 0 67068 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_89_730
timestamp 1562078211
transform 1 0 68172 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_89_742
timestamp 1562078211
transform 1 0 69276 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_754
timestamp 1
transform 1 0 70380 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_89_757
timestamp 1562078211
transform 1 0 70656 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_89_769
timestamp 1562078211
transform 1 0 71760 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_89_781
timestamp 1562078211
transform 1 0 72864 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_89_793
timestamp 1
transform 1 0 73968 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_90_706
timestamp 1562078211
transform 1 0 65964 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_90_718
timestamp 1
transform 1 0 67068 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_726
timestamp 1
transform 1 0 67804 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_40_12  FILLER_90_729
timestamp 1562078211
transform 1 0 68080 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_90_741
timestamp 1562078211
transform 1 0 69184 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_90_753
timestamp 1562078211
transform 1 0 70288 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_90_765
timestamp 1562078211
transform 1 0 71392 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_90_777
timestamp 1
transform 1 0 72496 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_781
timestamp 1
transform 1 0 72864 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_783
timestamp 1
transform 1 0 73048 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_90_785
timestamp 1562078211
transform 1 0 73232 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_90_797
timestamp 1
transform 1 0 74336 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_91_703
timestamp 1562078211
transform 1 0 65688 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_91_715
timestamp 1562078211
transform 1 0 66792 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_91_727
timestamp 1562078211
transform 1 0 67896 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_91_739
timestamp 1562078211
transform 1 0 69000 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_91_751
timestamp 1
transform 1 0 70104 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_755
timestamp 1
transform 1 0 70472 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_91_757
timestamp 1562078211
transform 1 0 70656 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_91_769
timestamp 1562078211
transform 1 0 71760 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_91_781
timestamp 1562078211
transform 1 0 72864 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_91_793
timestamp 1
transform 1 0 73968 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_92_703
timestamp 1562078211
transform 1 0 65688 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_92_715
timestamp 1562078211
transform 1 0 66792 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_727
timestamp 1
transform 1 0 67896 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_92_729
timestamp 1562078211
transform 1 0 68080 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_92_741
timestamp 1562078211
transform 1 0 69184 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_92_753
timestamp 1562078211
transform 1 0 70288 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_92_765
timestamp 1562078211
transform 1 0 71392 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_92_777
timestamp 1
transform 1 0 72496 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_781
timestamp 1
transform 1 0 72864 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_783
timestamp 1
transform 1 0 73048 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_92_785
timestamp 1562078211
transform 1 0 73232 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_92_797
timestamp 1
transform 1 0 74336 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_93_703
timestamp 1562078211
transform 1 0 65688 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_93_715
timestamp 1562078211
transform 1 0 66792 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_93_727
timestamp 1562078211
transform 1 0 67896 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_93_739
timestamp 1562078211
transform 1 0 69000 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_93_751
timestamp 1
transform 1 0 70104 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_755
timestamp 1
transform 1 0 70472 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_93_757
timestamp 1562078211
transform 1 0 70656 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_93_769
timestamp 1562078211
transform 1 0 71760 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_93_781
timestamp 1562078211
transform 1 0 72864 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_93_793
timestamp 1
transform 1 0 73968 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_94_709
timestamp 1562078211
transform 1 0 66240 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_94_721
timestamp 1
transform 1 0 67344 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_725
timestamp 1
transform 1 0 67712 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_727
timestamp 1
transform 1 0 67896 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_94_729
timestamp 1562078211
transform 1 0 68080 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_94_741
timestamp 1562078211
transform 1 0 69184 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_94_753
timestamp 1562078211
transform 1 0 70288 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_94_765
timestamp 1562078211
transform 1 0 71392 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_94_777
timestamp 1
transform 1 0 72496 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_781
timestamp 1
transform 1 0 72864 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_783
timestamp 1
transform 1 0 73048 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_94_785
timestamp 1562078211
transform 1 0 73232 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_94_797
timestamp 1
transform 1 0 74336 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_95_703
timestamp 1562078211
transform 1 0 65688 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_95_715
timestamp 1562078211
transform 1 0 66792 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_95_727
timestamp 1562078211
transform 1 0 67896 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_95_739
timestamp 1562078211
transform 1 0 69000 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_95_751
timestamp 1
transform 1 0 70104 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_755
timestamp 1
transform 1 0 70472 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_95_757
timestamp 1562078211
transform 1 0 70656 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_95_769
timestamp 1562078211
transform 1 0 71760 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_95_781
timestamp 1562078211
transform 1 0 72864 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_95_793
timestamp 1
transform 1 0 73968 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_96_703
timestamp 1562078211
transform 1 0 65688 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_96_715
timestamp 1562078211
transform 1 0 66792 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_727
timestamp 1
transform 1 0 67896 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_96_729
timestamp 1562078211
transform 1 0 68080 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_96_741
timestamp 1562078211
transform 1 0 69184 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_96_753
timestamp 1562078211
transform 1 0 70288 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_96_765
timestamp 1562078211
transform 1 0 71392 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_96_777
timestamp 1
transform 1 0 72496 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_781
timestamp 1
transform 1 0 72864 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_96_783
timestamp 1
transform 1 0 73048 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_96_785
timestamp 1562078211
transform 1 0 73232 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_96_797
timestamp 1
transform 1 0 74336 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_97_703
timestamp 1562078211
transform 1 0 65688 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_97_715
timestamp 1562078211
transform 1 0 66792 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_97_727
timestamp 1562078211
transform 1 0 67896 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_97_739
timestamp 1562078211
transform 1 0 69000 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_97_751
timestamp 1
transform 1 0 70104 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_755
timestamp 1
transform 1 0 70472 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_97_757
timestamp 1562078211
transform 1 0 70656 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_97_769
timestamp 1562078211
transform 1 0 71760 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_97_781
timestamp 1562078211
transform 1 0 72864 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_97_793
timestamp 1
transform 1 0 73968 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_98_703
timestamp 1562078211
transform 1 0 65688 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_98_715
timestamp 1562078211
transform 1 0 66792 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_727
timestamp 1
transform 1 0 67896 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_98_729
timestamp 1562078211
transform 1 0 68080 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_98_741
timestamp 1562078211
transform 1 0 69184 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_98_753
timestamp 1562078211
transform 1 0 70288 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_98_765
timestamp 1562078211
transform 1 0 71392 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_98_777
timestamp 1
transform 1 0 72496 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_781
timestamp 1
transform 1 0 72864 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_98_783
timestamp 1
transform 1 0 73048 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_98_785
timestamp 1562078211
transform 1 0 73232 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_98_797
timestamp 1
transform 1 0 74336 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_99_703
timestamp 1562078211
transform 1 0 65688 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_99_715
timestamp 1562078211
transform 1 0 66792 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_99_727
timestamp 1562078211
transform 1 0 67896 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_99_739
timestamp 1562078211
transform 1 0 69000 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_99_751
timestamp 1
transform 1 0 70104 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_755
timestamp 1
transform 1 0 70472 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_99_757
timestamp 1562078211
transform 1 0 70656 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_99_769
timestamp 1562078211
transform 1 0 71760 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_99_781
timestamp 1562078211
transform 1 0 72864 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_99_793
timestamp 1
transform 1 0 73968 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_100_703
timestamp 1562078211
transform 1 0 65688 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_100_715
timestamp 1562078211
transform 1 0 66792 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_727
timestamp 1
transform 1 0 67896 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_100_729
timestamp 1562078211
transform 1 0 68080 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_100_741
timestamp 1562078211
transform 1 0 69184 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_100_753
timestamp 1562078211
transform 1 0 70288 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_100_765
timestamp 1562078211
transform 1 0 71392 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_100_777
timestamp 1
transform 1 0 72496 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_781
timestamp 1
transform 1 0 72864 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_783
timestamp 1
transform 1 0 73048 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_100_785
timestamp 1562078211
transform 1 0 73232 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_100_797
timestamp 1
transform 1 0 74336 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_101_703
timestamp 1562078211
transform 1 0 65688 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_101_715
timestamp 1562078211
transform 1 0 66792 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_101_727
timestamp 1562078211
transform 1 0 67896 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_101_739
timestamp 1562078211
transform 1 0 69000 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_101_751
timestamp 1
transform 1 0 70104 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_755
timestamp 1
transform 1 0 70472 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_101_757
timestamp 1562078211
transform 1 0 70656 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_101_769
timestamp 1562078211
transform 1 0 71760 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_101_781
timestamp 1562078211
transform 1 0 72864 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_101_793
timestamp 1
transform 1 0 73968 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_102_703
timestamp 1562078211
transform 1 0 65688 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_102_715
timestamp 1562078211
transform 1 0 66792 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_727
timestamp 1
transform 1 0 67896 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_102_729
timestamp 1562078211
transform 1 0 68080 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_102_741
timestamp 1562078211
transform 1 0 69184 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_102_753
timestamp 1562078211
transform 1 0 70288 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_102_765
timestamp 1562078211
transform 1 0 71392 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_102_777
timestamp 1
transform 1 0 72496 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_102_781
timestamp 1
transform 1 0 72864 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_102_783
timestamp 1
transform 1 0 73048 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_102_785
timestamp 1562078211
transform 1 0 73232 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_102_797
timestamp 1
transform 1 0 74336 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_103_703
timestamp 1562078211
transform 1 0 65688 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_103_715
timestamp 1562078211
transform 1 0 66792 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_103_727
timestamp 1562078211
transform 1 0 67896 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_103_739
timestamp 1562078211
transform 1 0 69000 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_103_751
timestamp 1
transform 1 0 70104 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_755
timestamp 1
transform 1 0 70472 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_103_757
timestamp 1562078211
transform 1 0 70656 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_103_769
timestamp 1562078211
transform 1 0 71760 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_103_781
timestamp 1562078211
transform 1 0 72864 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_103_793
timestamp 1
transform 1 0 73968 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_104_703
timestamp 1562078211
transform 1 0 65688 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_104_715
timestamp 1562078211
transform 1 0 66792 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_727
timestamp 1
transform 1 0 67896 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_104_729
timestamp 1562078211
transform 1 0 68080 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_104_741
timestamp 1562078211
transform 1 0 69184 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_104_753
timestamp 1562078211
transform 1 0 70288 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_104_765
timestamp 1562078211
transform 1 0 71392 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_104_777
timestamp 1
transform 1 0 72496 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_781
timestamp 1
transform 1 0 72864 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_104_783
timestamp 1
transform 1 0 73048 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_104_785
timestamp 1562078211
transform 1 0 73232 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_104_797
timestamp 1
transform 1 0 74336 0 1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_105_703
timestamp 1562078211
transform 1 0 65688 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_105_715
timestamp 1562078211
transform 1 0 66792 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_105_727
timestamp 1562078211
transform 1 0 67896 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_105_739
timestamp 1562078211
transform 1 0 69000 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_105_751
timestamp 1
transform 1 0 70104 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_755
timestamp 1
transform 1 0 70472 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_105_757
timestamp 1562078211
transform 1 0 70656 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_105_769
timestamp 1562078211
transform 1 0 71760 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_105_781
timestamp 1562078211
transform 1 0 72864 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_105_793
timestamp 1
transform 1 0 73968 0 -1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_106_703
timestamp 1562078211
transform 1 0 65688 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_106_715
timestamp 1562078211
transform 1 0 66792 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_727
timestamp 1
transform 1 0 67896 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_106_729
timestamp 1562078211
transform 1 0 68080 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_106_741
timestamp 1562078211
transform 1 0 69184 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_106_753
timestamp 1562078211
transform 1 0 70288 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_106_765
timestamp 1562078211
transform 1 0 71392 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_106_777
timestamp 1
transform 1 0 72496 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_781
timestamp 1
transform 1 0 72864 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_106_783
timestamp 1
transform 1 0 73048 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_106_785
timestamp 1562078211
transform 1 0 73232 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_106_797
timestamp 1
transform 1 0 74336 0 1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_107_703
timestamp 1562078211
transform 1 0 65688 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_107_715
timestamp 1562078211
transform 1 0 66792 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_107_727
timestamp 1562078211
transform 1 0 67896 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_107_739
timestamp 1562078211
transform 1 0 69000 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_107_751
timestamp 1
transform 1 0 70104 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_755
timestamp 1
transform 1 0 70472 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_107_757
timestamp 1562078211
transform 1 0 70656 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_107_769
timestamp 1562078211
transform 1 0 71760 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_107_781
timestamp 1562078211
transform 1 0 72864 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_107_793
timestamp 1
transform 1 0 73968 0 -1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_108_703
timestamp 1562078211
transform 1 0 65688 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_108_715
timestamp 1562078211
transform 1 0 66792 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_727
timestamp 1
transform 1 0 67896 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_108_729
timestamp 1562078211
transform 1 0 68080 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_108_741
timestamp 1562078211
transform 1 0 69184 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_108_753
timestamp 1562078211
transform 1 0 70288 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_108_765
timestamp 1562078211
transform 1 0 71392 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_108_777
timestamp 1
transform 1 0 72496 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_781
timestamp 1
transform 1 0 72864 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_108_783
timestamp 1
transform 1 0 73048 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_108_785
timestamp 1562078211
transform 1 0 73232 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_108_797
timestamp 1
transform 1 0 74336 0 1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_109_703
timestamp 1562078211
transform 1 0 65688 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_109_715
timestamp 1562078211
transform 1 0 66792 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_109_727
timestamp 1562078211
transform 1 0 67896 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_109_739
timestamp 1562078211
transform 1 0 69000 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_109_751
timestamp 1
transform 1 0 70104 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_755
timestamp 1
transform 1 0 70472 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_109_757
timestamp 1562078211
transform 1 0 70656 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_109_769
timestamp 1562078211
transform 1 0 71760 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_109_781
timestamp 1562078211
transform 1 0 72864 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_109_793
timestamp 1
transform 1 0 73968 0 -1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_110_703
timestamp 1562078211
transform 1 0 65688 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_110_715
timestamp 1562078211
transform 1 0 66792 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_727
timestamp 1
transform 1 0 67896 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_110_729
timestamp 1562078211
transform 1 0 68080 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_110_741
timestamp 1562078211
transform 1 0 69184 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_110_753
timestamp 1562078211
transform 1 0 70288 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_110_765
timestamp 1562078211
transform 1 0 71392 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_110_777
timestamp 1
transform 1 0 72496 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_110_781
timestamp 1
transform 1 0 72864 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_110_783
timestamp 1
transform 1 0 73048 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_110_785
timestamp 1562078211
transform 1 0 73232 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_110_797
timestamp 1
transform 1 0 74336 0 1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_111_703
timestamp 1562078211
transform 1 0 65688 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_111_715
timestamp 1562078211
transform 1 0 66792 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_111_727
timestamp 1562078211
transform 1 0 67896 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_111_739
timestamp 1562078211
transform 1 0 69000 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_111_751
timestamp 1
transform 1 0 70104 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_755
timestamp 1
transform 1 0 70472 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_111_757
timestamp 1562078211
transform 1 0 70656 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_111_769
timestamp 1562078211
transform 1 0 71760 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_111_781
timestamp 1562078211
transform 1 0 72864 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_111_793
timestamp 1
transform 1 0 73968 0 -1 62016
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_112_703
timestamp 1562078211
transform 1 0 65688 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_112_715
timestamp 1562078211
transform 1 0 66792 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_727
timestamp 1
transform 1 0 67896 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_112_729
timestamp 1562078211
transform 1 0 68080 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_112_741
timestamp 1562078211
transform 1 0 69184 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_112_753
timestamp 1562078211
transform 1 0 70288 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_112_765
timestamp 1562078211
transform 1 0 71392 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_112_777
timestamp 1
transform 1 0 72496 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_112_781
timestamp 1
transform 1 0 72864 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_112_783
timestamp 1
transform 1 0 73048 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_112_785
timestamp 1562078211
transform 1 0 73232 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_112_797
timestamp 1
transform 1 0 74336 0 1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_113_703
timestamp 1562078211
transform 1 0 65688 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_113_715
timestamp 1562078211
transform 1 0 66792 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_113_727
timestamp 1562078211
transform 1 0 67896 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_113_739
timestamp 1562078211
transform 1 0 69000 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_113_751
timestamp 1
transform 1 0 70104 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_755
timestamp 1
transform 1 0 70472 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_113_757
timestamp 1562078211
transform 1 0 70656 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_113_769
timestamp 1562078211
transform 1 0 71760 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_113_781
timestamp 1562078211
transform 1 0 72864 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_113_793
timestamp 1
transform 1 0 73968 0 -1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_114_703
timestamp 1562078211
transform 1 0 65688 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_114_715
timestamp 1562078211
transform 1 0 66792 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_727
timestamp 1
transform 1 0 67896 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_114_729
timestamp 1562078211
transform 1 0 68080 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_114_741
timestamp 1562078211
transform 1 0 69184 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_114_753
timestamp 1562078211
transform 1 0 70288 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_114_765
timestamp 1562078211
transform 1 0 71392 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_114_777
timestamp 1
transform 1 0 72496 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_114_781
timestamp 1
transform 1 0 72864 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_114_783
timestamp 1
transform 1 0 73048 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_114_785
timestamp 1562078211
transform 1 0 73232 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_114_797
timestamp 1
transform 1 0 74336 0 1 63104
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_115_703
timestamp 1562078211
transform 1 0 65688 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_115_715
timestamp 1562078211
transform 1 0 66792 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_115_727
timestamp 1562078211
transform 1 0 67896 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_115_739
timestamp 1562078211
transform 1 0 69000 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_115_751
timestamp 1
transform 1 0 70104 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_755
timestamp 1
transform 1 0 70472 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_115_757
timestamp 1562078211
transform 1 0 70656 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_115_769
timestamp 1562078211
transform 1 0 71760 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_115_781
timestamp 1562078211
transform 1 0 72864 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_115_793
timestamp 1
transform 1 0 73968 0 -1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_116_703
timestamp 1562078211
transform 1 0 65688 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_116_715
timestamp 1562078211
transform 1 0 66792 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_727
timestamp 1
transform 1 0 67896 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_116_729
timestamp 1562078211
transform 1 0 68080 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_116_741
timestamp 1562078211
transform 1 0 69184 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_116_753
timestamp 1562078211
transform 1 0 70288 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_116_765
timestamp 1562078211
transform 1 0 71392 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_116_777
timestamp 1
transform 1 0 72496 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_116_781
timestamp 1
transform 1 0 72864 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_116_783
timestamp 1
transform 1 0 73048 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_116_785
timestamp 1562078211
transform 1 0 73232 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_116_797
timestamp 1
transform 1 0 74336 0 1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_117_703
timestamp 1562078211
transform 1 0 65688 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_117_715
timestamp 1562078211
transform 1 0 66792 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_117_727
timestamp 1562078211
transform 1 0 67896 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_117_739
timestamp 1562078211
transform 1 0 69000 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_117_751
timestamp 1
transform 1 0 70104 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_755
timestamp 1
transform 1 0 70472 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_117_757
timestamp 1562078211
transform 1 0 70656 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_117_769
timestamp 1562078211
transform 1 0 71760 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_117_781
timestamp 1562078211
transform 1 0 72864 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_117_793
timestamp 1
transform 1 0 73968 0 -1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_118_703
timestamp 1562078211
transform 1 0 65688 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_118_715
timestamp 1562078211
transform 1 0 66792 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_727
timestamp 1
transform 1 0 67896 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_118_729
timestamp 1562078211
transform 1 0 68080 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_118_741
timestamp 1562078211
transform 1 0 69184 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_118_753
timestamp 1562078211
transform 1 0 70288 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_118_765
timestamp 1562078211
transform 1 0 71392 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_118_777
timestamp 1
transform 1 0 72496 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_118_781
timestamp 1
transform 1 0 72864 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_118_783
timestamp 1
transform 1 0 73048 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_118_785
timestamp 1562078211
transform 1 0 73232 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_118_797
timestamp 1
transform 1 0 74336 0 1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_119_703
timestamp 1562078211
transform 1 0 65688 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_119_715
timestamp 1562078211
transform 1 0 66792 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_119_727
timestamp 1562078211
transform 1 0 67896 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_119_739
timestamp 1562078211
transform 1 0 69000 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_119_751
timestamp 1
transform 1 0 70104 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_755
timestamp 1
transform 1 0 70472 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_119_757
timestamp 1562078211
transform 1 0 70656 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_119_769
timestamp 1562078211
transform 1 0 71760 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_119_781
timestamp 1562078211
transform 1 0 72864 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_119_793
timestamp 1
transform 1 0 73968 0 -1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_120_703
timestamp 1562078211
transform 1 0 65688 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_120_715
timestamp 1562078211
transform 1 0 66792 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_727
timestamp 1
transform 1 0 67896 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_120_729
timestamp 1562078211
transform 1 0 68080 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_120_741
timestamp 1562078211
transform 1 0 69184 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_120_753
timestamp 1562078211
transform 1 0 70288 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_120_765
timestamp 1562078211
transform 1 0 71392 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_120_777
timestamp 1
transform 1 0 72496 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_120_781
timestamp 1
transform 1 0 72864 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_120_783
timestamp 1
transform 1 0 73048 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_120_785
timestamp 1562078211
transform 1 0 73232 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_120_797
timestamp 1
transform 1 0 74336 0 1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_121_703
timestamp 1562078211
transform 1 0 65688 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_121_715
timestamp 1562078211
transform 1 0 66792 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_121_727
timestamp 1562078211
transform 1 0 67896 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_121_739
timestamp 1562078211
transform 1 0 69000 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_121_751
timestamp 1
transform 1 0 70104 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_755
timestamp 1
transform 1 0 70472 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_121_757
timestamp 1562078211
transform 1 0 70656 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_121_769
timestamp 1562078211
transform 1 0 71760 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_121_781
timestamp 1562078211
transform 1 0 72864 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_121_793
timestamp 1
transform 1 0 73968 0 -1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_122_703
timestamp 1562078211
transform 1 0 65688 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_122_715
timestamp 1562078211
transform 1 0 66792 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_727
timestamp 1
transform 1 0 67896 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_122_729
timestamp 1562078211
transform 1 0 68080 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_122_741
timestamp 1562078211
transform 1 0 69184 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_122_753
timestamp 1562078211
transform 1 0 70288 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_122_765
timestamp 1562078211
transform 1 0 71392 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_122_777
timestamp 1
transform 1 0 72496 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_122_781
timestamp 1
transform 1 0 72864 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_122_783
timestamp 1
transform 1 0 73048 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_122_785
timestamp 1562078211
transform 1 0 73232 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_122_797
timestamp 1
transform 1 0 74336 0 1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_123_703
timestamp 1562078211
transform 1 0 65688 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_123_715
timestamp 1562078211
transform 1 0 66792 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_123_727
timestamp 1562078211
transform 1 0 67896 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_123_739
timestamp 1562078211
transform 1 0 69000 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_123_751
timestamp 1
transform 1 0 70104 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_755
timestamp 1
transform 1 0 70472 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_123_757
timestamp 1562078211
transform 1 0 70656 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_123_769
timestamp 1562078211
transform 1 0 71760 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_123_781
timestamp 1562078211
transform 1 0 72864 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_123_793
timestamp 1
transform 1 0 73968 0 -1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_124_703
timestamp 1562078211
transform 1 0 65688 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_124_715
timestamp 1562078211
transform 1 0 66792 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_727
timestamp 1
transform 1 0 67896 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_124_729
timestamp 1562078211
transform 1 0 68080 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_124_741
timestamp 1562078211
transform 1 0 69184 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_124_753
timestamp 1562078211
transform 1 0 70288 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_124_765
timestamp 1562078211
transform 1 0 71392 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_124_777
timestamp 1
transform 1 0 72496 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_124_781
timestamp 1
transform 1 0 72864 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_124_783
timestamp 1
transform 1 0 73048 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_124_785
timestamp 1562078211
transform 1 0 73232 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_124_797
timestamp 1
transform 1 0 74336 0 1 68544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_125_703
timestamp 1562078211
transform 1 0 65688 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_125_715
timestamp 1562078211
transform 1 0 66792 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_125_727
timestamp 1562078211
transform 1 0 67896 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_125_739
timestamp 1562078211
transform 1 0 69000 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_125_751
timestamp 1
transform 1 0 70104 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_755
timestamp 1
transform 1 0 70472 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_125_757
timestamp 1562078211
transform 1 0 70656 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_125_769
timestamp 1562078211
transform 1 0 71760 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_125_781
timestamp 1562078211
transform 1 0 72864 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_125_793
timestamp 1
transform 1 0 73968 0 -1 69632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_126_703
timestamp 1562078211
transform 1 0 65688 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_126_715
timestamp 1562078211
transform 1 0 66792 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_727
timestamp 1
transform 1 0 67896 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_126_729
timestamp 1562078211
transform 1 0 68080 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_126_741
timestamp 1562078211
transform 1 0 69184 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_126_753
timestamp 1562078211
transform 1 0 70288 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_126_765
timestamp 1562078211
transform 1 0 71392 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_126_777
timestamp 1
transform 1 0 72496 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_126_781
timestamp 1
transform 1 0 72864 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_126_783
timestamp 1
transform 1 0 73048 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_126_785
timestamp 1562078211
transform 1 0 73232 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_126_797
timestamp 1
transform 1 0 74336 0 1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_127_703
timestamp 1562078211
transform 1 0 65688 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_127_715
timestamp 1562078211
transform 1 0 66792 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_127_727
timestamp 1562078211
transform 1 0 67896 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_127_739
timestamp 1562078211
transform 1 0 69000 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_127_751
timestamp 1
transform 1 0 70104 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_755
timestamp 1
transform 1 0 70472 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_127_757
timestamp 1562078211
transform 1 0 70656 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_127_769
timestamp 1562078211
transform 1 0 71760 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_127_781
timestamp 1562078211
transform 1 0 72864 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_127_793
timestamp 1
transform 1 0 73968 0 -1 70720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_128_703
timestamp 1562078211
transform 1 0 65688 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_128_715
timestamp 1562078211
transform 1 0 66792 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_727
timestamp 1
transform 1 0 67896 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_128_729
timestamp 1562078211
transform 1 0 68080 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_128_741
timestamp 1562078211
transform 1 0 69184 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_128_753
timestamp 1562078211
transform 1 0 70288 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_128_765
timestamp 1562078211
transform 1 0 71392 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_128_777
timestamp 1
transform 1 0 72496 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_128_781
timestamp 1
transform 1 0 72864 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_128_783
timestamp 1
transform 1 0 73048 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_128_785
timestamp 1562078211
transform 1 0 73232 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_128_797
timestamp 1
transform 1 0 74336 0 1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_129_703
timestamp 1562078211
transform 1 0 65688 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_129_715
timestamp 1562078211
transform 1 0 66792 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_129_727
timestamp 1562078211
transform 1 0 67896 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_129_739
timestamp 1562078211
transform 1 0 69000 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_129_751
timestamp 1
transform 1 0 70104 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_755
timestamp 1
transform 1 0 70472 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_129_757
timestamp 1562078211
transform 1 0 70656 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_129_769
timestamp 1562078211
transform 1 0 71760 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_129_781
timestamp 1562078211
transform 1 0 72864 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_129_793
timestamp 1
transform 1 0 73968 0 -1 71808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_130_703
timestamp 1562078211
transform 1 0 65688 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_130_715
timestamp 1562078211
transform 1 0 66792 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_727
timestamp 1
transform 1 0 67896 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_130_729
timestamp 1562078211
transform 1 0 68080 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_130_741
timestamp 1562078211
transform 1 0 69184 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_130_753
timestamp 1562078211
transform 1 0 70288 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_130_765
timestamp 1562078211
transform 1 0 71392 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_130_777
timestamp 1
transform 1 0 72496 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_130_781
timestamp 1
transform 1 0 72864 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_130_783
timestamp 1
transform 1 0 73048 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_130_785
timestamp 1562078211
transform 1 0 73232 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_130_797
timestamp 1
transform 1 0 74336 0 1 71808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_131_703
timestamp 1562078211
transform 1 0 65688 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_131_715
timestamp 1562078211
transform 1 0 66792 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_131_727
timestamp 1562078211
transform 1 0 67896 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_131_739
timestamp 1562078211
transform 1 0 69000 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_131_751
timestamp 1
transform 1 0 70104 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_755
timestamp 1
transform 1 0 70472 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_131_757
timestamp 1562078211
transform 1 0 70656 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_131_769
timestamp 1562078211
transform 1 0 71760 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_131_781
timestamp 1562078211
transform 1 0 72864 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_131_793
timestamp 1
transform 1 0 73968 0 -1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_132_703
timestamp 1562078211
transform 1 0 65688 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_132_715
timestamp 1562078211
transform 1 0 66792 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_727
timestamp 1
transform 1 0 67896 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_132_729
timestamp 1562078211
transform 1 0 68080 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_132_741
timestamp 1562078211
transform 1 0 69184 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_132_753
timestamp 1562078211
transform 1 0 70288 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_132_765
timestamp 1562078211
transform 1 0 71392 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_132_777
timestamp 1
transform 1 0 72496 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_132_781
timestamp 1
transform 1 0 72864 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_132_783
timestamp 1
transform 1 0 73048 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_132_785
timestamp 1562078211
transform 1 0 73232 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_132_797
timestamp 1
transform 1 0 74336 0 1 72896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_133_703
timestamp 1562078211
transform 1 0 65688 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_133_715
timestamp 1562078211
transform 1 0 66792 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_133_727
timestamp 1562078211
transform 1 0 67896 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_133_739
timestamp 1562078211
transform 1 0 69000 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_133_751
timestamp 1
transform 1 0 70104 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_755
timestamp 1
transform 1 0 70472 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_133_757
timestamp 1562078211
transform 1 0 70656 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_133_769
timestamp 1562078211
transform 1 0 71760 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_133_781
timestamp 1562078211
transform 1 0 72864 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_133_793
timestamp 1
transform 1 0 73968 0 -1 73984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_134_703
timestamp 1562078211
transform 1 0 65688 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_134_715
timestamp 1562078211
transform 1 0 66792 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_727
timestamp 1
transform 1 0 67896 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_134_729
timestamp 1562078211
transform 1 0 68080 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_134_741
timestamp 1562078211
transform 1 0 69184 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_134_753
timestamp 1562078211
transform 1 0 70288 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_134_765
timestamp 1562078211
transform 1 0 71392 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_134_777
timestamp 1
transform 1 0 72496 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_134_781
timestamp 1
transform 1 0 72864 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_134_783
timestamp 1
transform 1 0 73048 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_134_785
timestamp 1562078211
transform 1 0 73232 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_134_797
timestamp 1
transform 1 0 74336 0 1 73984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_135_703
timestamp 1562078211
transform 1 0 65688 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_135_715
timestamp 1562078211
transform 1 0 66792 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_135_727
timestamp 1562078211
transform 1 0 67896 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_135_739
timestamp 1562078211
transform 1 0 69000 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_135_751
timestamp 1
transform 1 0 70104 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_755
timestamp 1
transform 1 0 70472 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_135_757
timestamp 1562078211
transform 1 0 70656 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_135_769
timestamp 1562078211
transform 1 0 71760 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_135_781
timestamp 1562078211
transform 1 0 72864 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_135_793
timestamp 1
transform 1 0 73968 0 -1 75072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_136_703
timestamp 1562078211
transform 1 0 65688 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_136_715
timestamp 1562078211
transform 1 0 66792 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_727
timestamp 1
transform 1 0 67896 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_136_729
timestamp 1562078211
transform 1 0 68080 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_136_741
timestamp 1562078211
transform 1 0 69184 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_136_753
timestamp 1562078211
transform 1 0 70288 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_136_765
timestamp 1562078211
transform 1 0 71392 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_136_777
timestamp 1
transform 1 0 72496 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_136_781
timestamp 1
transform 1 0 72864 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_136_783
timestamp 1
transform 1 0 73048 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_136_785
timestamp 1562078211
transform 1 0 73232 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_136_797
timestamp 1
transform 1 0 74336 0 1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_137_703
timestamp 1562078211
transform 1 0 65688 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_137_715
timestamp 1562078211
transform 1 0 66792 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_137_727
timestamp 1562078211
transform 1 0 67896 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_137_739
timestamp 1562078211
transform 1 0 69000 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_137_751
timestamp 1
transform 1 0 70104 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_755
timestamp 1
transform 1 0 70472 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_137_757
timestamp 1562078211
transform 1 0 70656 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_137_769
timestamp 1562078211
transform 1 0 71760 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_137_781
timestamp 1562078211
transform 1 0 72864 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_137_793
timestamp 1
transform 1 0 73968 0 -1 76160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_138_703
timestamp 1562078211
transform 1 0 65688 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_138_715
timestamp 1562078211
transform 1 0 66792 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_727
timestamp 1
transform 1 0 67896 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_138_729
timestamp 1562078211
transform 1 0 68080 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_138_741
timestamp 1562078211
transform 1 0 69184 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_138_753
timestamp 1562078211
transform 1 0 70288 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_138_765
timestamp 1562078211
transform 1 0 71392 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_138_777
timestamp 1
transform 1 0 72496 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_138_781
timestamp 1
transform 1 0 72864 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_138_783
timestamp 1
transform 1 0 73048 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_138_785
timestamp 1562078211
transform 1 0 73232 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_138_797
timestamp 1
transform 1 0 74336 0 1 76160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_139_703
timestamp 1562078211
transform 1 0 65688 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_139_715
timestamp 1562078211
transform 1 0 66792 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_139_727
timestamp 1562078211
transform 1 0 67896 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_139_739
timestamp 1562078211
transform 1 0 69000 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_139_751
timestamp 1
transform 1 0 70104 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_139_755
timestamp 1
transform 1 0 70472 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_139_757
timestamp 1562078211
transform 1 0 70656 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_139_769
timestamp 1562078211
transform 1 0 71760 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_139_781
timestamp 1562078211
transform 1 0 72864 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_139_793
timestamp 1
transform 1 0 73968 0 -1 77248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_140_703
timestamp 1562078211
transform 1 0 65688 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_140_715
timestamp 1562078211
transform 1 0 66792 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_727
timestamp 1
transform 1 0 67896 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_140_729
timestamp 1562078211
transform 1 0 68080 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_140_741
timestamp 1562078211
transform 1 0 69184 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_140_753
timestamp 1562078211
transform 1 0 70288 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_140_765
timestamp 1562078211
transform 1 0 71392 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_140_777
timestamp 1
transform 1 0 72496 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_140_781
timestamp 1
transform 1 0 72864 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_140_783
timestamp 1
transform 1 0 73048 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_140_785
timestamp 1562078211
transform 1 0 73232 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_140_797
timestamp 1
transform 1 0 74336 0 1 77248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_141_703
timestamp 1562078211
transform 1 0 65688 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_141_715
timestamp 1562078211
transform 1 0 66792 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_141_727
timestamp 1562078211
transform 1 0 67896 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_141_739
timestamp 1562078211
transform 1 0 69000 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_141_751
timestamp 1
transform 1 0 70104 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_141_755
timestamp 1
transform 1 0 70472 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_141_757
timestamp 1562078211
transform 1 0 70656 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_141_769
timestamp 1562078211
transform 1 0 71760 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_141_781
timestamp 1562078211
transform 1 0 72864 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_141_793
timestamp 1
transform 1 0 73968 0 -1 78336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_142_703
timestamp 1562078211
transform 1 0 65688 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_142_715
timestamp 1562078211
transform 1 0 66792 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_727
timestamp 1
transform 1 0 67896 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_142_729
timestamp 1562078211
transform 1 0 68080 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_142_741
timestamp 1562078211
transform 1 0 69184 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_142_753
timestamp 1562078211
transform 1 0 70288 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_142_765
timestamp 1562078211
transform 1 0 71392 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_142_777
timestamp 1
transform 1 0 72496 0 1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_142_781
timestamp 1
transform 1 0 72864 0 1 78336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_142_783
timestamp 1
transform 1 0 73048 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_142_785
timestamp 1562078211
transform 1 0 73232 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_142_797
timestamp 1
transform 1 0 74336 0 1 78336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_143_703
timestamp 1562078211
transform 1 0 65688 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_143_715
timestamp 1562078211
transform 1 0 66792 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_143_727
timestamp 1562078211
transform 1 0 67896 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_143_739
timestamp 1562078211
transform 1 0 69000 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_143_751
timestamp 1
transform 1 0 70104 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_143_755
timestamp 1
transform 1 0 70472 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_143_757
timestamp 1562078211
transform 1 0 70656 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_143_769
timestamp 1562078211
transform 1 0 71760 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_143_781
timestamp 1562078211
transform 1 0 72864 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_143_793
timestamp 1
transform 1 0 73968 0 -1 79424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_144_703
timestamp 1562078211
transform 1 0 65688 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_144_715
timestamp 1562078211
transform 1 0 66792 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_727
timestamp 1
transform 1 0 67896 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_144_729
timestamp 1562078211
transform 1 0 68080 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_144_741
timestamp 1562078211
transform 1 0 69184 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_144_753
timestamp 1562078211
transform 1 0 70288 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_144_765
timestamp 1562078211
transform 1 0 71392 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_144_777
timestamp 1
transform 1 0 72496 0 1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_144_781
timestamp 1
transform 1 0 72864 0 1 79424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_144_783
timestamp 1
transform 1 0 73048 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_144_785
timestamp 1562078211
transform 1 0 73232 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_144_797
timestamp 1
transform 1 0 74336 0 1 79424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_145_703
timestamp 1562078211
transform 1 0 65688 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_145_715
timestamp 1562078211
transform 1 0 66792 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_145_727
timestamp 1562078211
transform 1 0 67896 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_145_739
timestamp 1562078211
transform 1 0 69000 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_145_751
timestamp 1
transform 1 0 70104 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_145_755
timestamp 1
transform 1 0 70472 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_145_757
timestamp 1562078211
transform 1 0 70656 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_145_769
timestamp 1562078211
transform 1 0 71760 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_145_781
timestamp 1562078211
transform 1 0 72864 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_145_793
timestamp 1
transform 1 0 73968 0 -1 80512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_146_703
timestamp 1562078211
transform 1 0 65688 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_146_715
timestamp 1562078211
transform 1 0 66792 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_727
timestamp 1
transform 1 0 67896 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_146_729
timestamp 1562078211
transform 1 0 68080 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_146_741
timestamp 1562078211
transform 1 0 69184 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_146_753
timestamp 1562078211
transform 1 0 70288 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_146_765
timestamp 1562078211
transform 1 0 71392 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_146_777
timestamp 1
transform 1 0 72496 0 1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_146_781
timestamp 1
transform 1 0 72864 0 1 80512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_146_783
timestamp 1
transform 1 0 73048 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_146_785
timestamp 1562078211
transform 1 0 73232 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_146_797
timestamp 1
transform 1 0 74336 0 1 80512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_147_703
timestamp 1562078211
transform 1 0 65688 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_147_715
timestamp 1562078211
transform 1 0 66792 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_147_727
timestamp 1562078211
transform 1 0 67896 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_147_739
timestamp 1562078211
transform 1 0 69000 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_147_751
timestamp 1
transform 1 0 70104 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_147_755
timestamp 1
transform 1 0 70472 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_147_757
timestamp 1562078211
transform 1 0 70656 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_147_769
timestamp 1562078211
transform 1 0 71760 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_147_781
timestamp 1562078211
transform 1 0 72864 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_147_793
timestamp 1
transform 1 0 73968 0 -1 81600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_148_703
timestamp 1562078211
transform 1 0 65688 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_148_715
timestamp 1562078211
transform 1 0 66792 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_727
timestamp 1
transform 1 0 67896 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_148_729
timestamp 1562078211
transform 1 0 68080 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_148_741
timestamp 1562078211
transform 1 0 69184 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_148_753
timestamp 1562078211
transform 1 0 70288 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_148_765
timestamp 1562078211
transform 1 0 71392 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_148_777
timestamp 1
transform 1 0 72496 0 1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_148_781
timestamp 1
transform 1 0 72864 0 1 81600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_148_783
timestamp 1
transform 1 0 73048 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_148_785
timestamp 1562078211
transform 1 0 73232 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_148_797
timestamp 1
transform 1 0 74336 0 1 81600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_149_703
timestamp 1562078211
transform 1 0 65688 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_149_715
timestamp 1562078211
transform 1 0 66792 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_149_727
timestamp 1562078211
transform 1 0 67896 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_149_739
timestamp 1562078211
transform 1 0 69000 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_149_751
timestamp 1
transform 1 0 70104 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_755
timestamp 1
transform 1 0 70472 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_149_757
timestamp 1562078211
transform 1 0 70656 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_149_769
timestamp 1562078211
transform 1 0 71760 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_149_781
timestamp 1562078211
transform 1 0 72864 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_149_793
timestamp 1
transform 1 0 73968 0 -1 82688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_150_703
timestamp 1562078211
transform 1 0 65688 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_150_715
timestamp 1562078211
transform 1 0 66792 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_727
timestamp 1
transform 1 0 67896 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_150_729
timestamp 1562078211
transform 1 0 68080 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_150_741
timestamp 1562078211
transform 1 0 69184 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_150_753
timestamp 1562078211
transform 1 0 70288 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_150_765
timestamp 1562078211
transform 1 0 71392 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_150_777
timestamp 1
transform 1 0 72496 0 1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_150_781
timestamp 1
transform 1 0 72864 0 1 82688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_150_783
timestamp 1
transform 1 0 73048 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_150_785
timestamp 1562078211
transform 1 0 73232 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_150_797
timestamp 1
transform 1 0 74336 0 1 82688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_151_703
timestamp 1562078211
transform 1 0 65688 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_151_715
timestamp 1562078211
transform 1 0 66792 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_151_727
timestamp 1562078211
transform 1 0 67896 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_151_739
timestamp 1562078211
transform 1 0 69000 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_151_751
timestamp 1
transform 1 0 70104 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_755
timestamp 1
transform 1 0 70472 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_151_757
timestamp 1562078211
transform 1 0 70656 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_151_769
timestamp 1562078211
transform 1 0 71760 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_151_781
timestamp 1562078211
transform 1 0 72864 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_151_793
timestamp 1
transform 1 0 73968 0 -1 83776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_152_703
timestamp 1562078211
transform 1 0 65688 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_152_715
timestamp 1562078211
transform 1 0 66792 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_727
timestamp 1
transform 1 0 67896 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_152_729
timestamp 1562078211
transform 1 0 68080 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_152_741
timestamp 1562078211
transform 1 0 69184 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_152_753
timestamp 1562078211
transform 1 0 70288 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_152_765
timestamp 1562078211
transform 1 0 71392 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_152_777
timestamp 1
transform 1 0 72496 0 1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_152_781
timestamp 1
transform 1 0 72864 0 1 83776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_152_783
timestamp 1
transform 1 0 73048 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_152_785
timestamp 1562078211
transform 1 0 73232 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_152_797
timestamp 1
transform 1 0 74336 0 1 83776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_153_703
timestamp 1562078211
transform 1 0 65688 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_153_715
timestamp 1562078211
transform 1 0 66792 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_153_727
timestamp 1562078211
transform 1 0 67896 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_153_739
timestamp 1562078211
transform 1 0 69000 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_153_751
timestamp 1
transform 1 0 70104 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_755
timestamp 1
transform 1 0 70472 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_153_757
timestamp 1562078211
transform 1 0 70656 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_153_769
timestamp 1562078211
transform 1 0 71760 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_153_781
timestamp 1562078211
transform 1 0 72864 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_8  FILLER_153_793
timestamp 1
transform 1 0 73968 0 -1 84864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_40_12  FILLER_154_703
timestamp 1562078211
transform 1 0 65688 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_154_715
timestamp 1562078211
transform 1 0 66792 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_727
timestamp 1
transform 1 0 67896 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_154_729
timestamp 1562078211
transform 1 0 68080 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_154_741
timestamp 1562078211
transform 1 0 69184 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_154_753
timestamp 1562078211
transform 1 0 70288 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_154_765
timestamp 1562078211
transform 1 0 71392 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_154_777
timestamp 1
transform 1 0 72496 0 1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_154_781
timestamp 1
transform 1 0 72864 0 1 84864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_154_783
timestamp 1
transform 1 0 73048 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_154_785
timestamp 1562078211
transform 1 0 73232 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_154_797
timestamp 1
transform 1 0 74336 0 1 84864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_40_12  FILLER_155_703
timestamp 1562078211
transform 1 0 65688 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_155_715
timestamp 1562078211
transform 1 0 66792 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_155_727
timestamp 1
transform 1 0 67896 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_155_729
timestamp 1562078211
transform 1 0 68080 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_155_741
timestamp 1562078211
transform 1 0 69184 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_155_753
timestamp 1
transform 1 0 70288 0 -1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_155_755
timestamp 1
transform 1 0 70472 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_155_757
timestamp 1562078211
transform 1 0 70656 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_40_12  FILLER_155_769
timestamp 1562078211
transform 1 0 71760 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_155_781
timestamp 1
transform 1 0 72864 0 -1 85952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_155_783
timestamp 1
transform 1 0 73048 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_40_12  FILLER_155_785
timestamp 1562078211
transform 1 0 73232 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_155_797
timestamp 1
transform 1 0 74336 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 49680 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 56672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform 1 0 27876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform 1 0 47472 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 43148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform 1 0 53360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform 1 0 66608 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 66424 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform 1 0 26036 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform 1 0 44068 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform 1 0 67068 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 66424 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform 1 0 40940 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform 1 0 52624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform 1 0 24564 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform 1 0 44804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 49680 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform 1 0 55936 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform 1 0 69368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 67160 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform 1 0 46368 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform 1 0 55200 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 39928 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform 1 0 51520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform 1 0 70656 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform -1 0 67436 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform 1 0 45080 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform 1 0 54280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 73968 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 68816 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform 1 0 37720 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform 1 0 50508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform 1 0 35604 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform 1 0 50784 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform 1 0 43884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform 1 0 54096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform 1 0 32200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform 1 0 50048 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform 1 0 53544 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform -1 0 66424 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform 1 0 43884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 67344 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform 1 0 51612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform -1 0 66424 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform 1 0 55200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform -1 0 66424 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform 1 0 32936 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform 1 0 48944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1
transform -1 0 52256 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1
transform -1 0 66424 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1
transform 1 0 56212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1
transform -1 0 66424 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1
transform -1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1
transform -1 0 66424 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1
transform -1 0 59984 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1
transform -1 0 66424 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1
transform -1 0 60168 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1
transform -1 0 66424 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1
transform -1 0 62008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1
transform -1 0 66424 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1
transform -1 0 41400 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1
transform -1 0 67896 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1
transform 1 0 62192 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1
transform -1 0 66424 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1
transform -1 0 30728 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1
transform 1 0 48392 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1
transform -1 0 67160 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1
transform 1 0 37076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1
transform -1 0 67344 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1
transform 1 0 31464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1
transform -1 0 66608 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1
transform 1 0 63664 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1
transform -1 0 66424 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1
transform 1 0 65504 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1
transform -1 0 66424 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1
transform 1 0 35972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1
transform -1 0 66424 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1
transform -1 0 66608 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1
transform -1 0 29348 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1
transform -1 0 66424 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1
transform -1 0 30268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1
transform -1 0 66792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1
transform 1 0 27324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold86
timestamp 1
transform 1 0 47472 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1
transform -1 0 29348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1
transform 1 0 27140 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold89
timestamp 1
transform 1 0 45540 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1
transform 1 0 28796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold92
timestamp 1
transform 1 0 65688 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1
transform 1 0 26036 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1
transform 1 0 32016 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold95
timestamp 1
transform 1 0 65688 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1
transform 1 0 27140 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1
transform -1 0 50140 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1
transform 1 0 47472 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1
transform 1 0 46276 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1
transform -1 0 47380 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1
transform -1 0 46092 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1
transform 1 0 42320 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1
transform -1 0 42136 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1
transform -1 0 40664 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1
transform -1 0 38548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1
transform 1 0 34776 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1
transform -1 0 54832 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1
transform -1 0 35788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1
transform -1 0 57408 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1
transform -1 0 53360 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1
transform 1 0 54924 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1
transform 1 0 59248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1
transform 1 0 50140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1
transform 1 0 57776 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1
transform -1 0 34408 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1
transform 1 0 60720 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1
transform 1 0 61272 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1
transform -1 0 28796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1
transform -1 0 31004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1
transform -1 0 66240 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1
transform 1 0 65688 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1
transform -1 0 28244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1
transform 1 0 66976 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1
transform 1 0 63848 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1
transform -1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1
transform -1 0 70288 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1
transform 1 0 68448 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1
transform 1 0 72128 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1
transform 1 0 43148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1
transform -1 0 44528 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1
transform -1 0 41952 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1
transform 1 0 37444 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1
transform 1 0 36340 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1
transform 1 0 29716 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1
transform -1 0 36708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1
transform 1 0 30728 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1
transform 1 0 25300 0 -1 2176
box -38 -48 774 592
use CF_SRAM_1024x32  i_sram
timestamp 1586029971
transform 0 -1 63375 1 0 8000
box 0 0 77574 61355
use sky130_fd_sc_hd__conb_1  i_sram_90
timestamp 1
transform -1 0 65964 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  i_sram_91
timestamp 1
transform -1 0 65964 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  i_sram_92
timestamp 1
transform -1 0 65964 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  i_sram_93
timestamp 1
transform -1 0 65964 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  i_sram_94
timestamp 1
transform -1 0 65964 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  i_sram_95
timestamp 1
transform -1 0 66240 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  i_sram_96
timestamp 1
transform -1 0 65964 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  i_sram_97
timestamp 1
transform 1 0 65688 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  i_sram_98
timestamp 1
transform 1 0 65964 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1
transform 1 0 23552 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1
transform -1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1
transform 1 0 44620 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input4
timestamp 1
transform -1 0 27140 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 1
transform -1 0 28980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input6
timestamp 1
transform -1 0 32844 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1
transform 1 0 35972 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1
transform -1 0 36432 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1
transform -1 0 37720 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1
transform -1 0 39192 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1
transform -1 0 40664 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1
transform 1 0 24196 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1
transform 1 0 25668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1
transform -1 0 42228 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1
transform 1 0 45172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1
transform 1 0 45816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1
transform 1 0 47012 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1
transform -1 0 47840 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1
transform -1 0 48944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1
transform -1 0 50692 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1
transform 1 0 52348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input22
timestamp 1
transform 1 0 54280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1
transform 1 0 55660 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input24
timestamp 1
transform -1 0 26772 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1
transform 1 0 56948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1
transform -1 0 58328 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input27
timestamp 1
transform -1 0 59800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input28
timestamp 1
transform -1 0 61272 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input29
timestamp 1
transform -1 0 62744 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1
transform 1 0 68080 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1
transform -1 0 66056 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input32
timestamp 1
transform 1 0 67344 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input33
timestamp 1
transform 1 0 68080 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input34
timestamp 1
transform 1 0 70840 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input35
timestamp 1
transform 1 0 29440 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input36
timestamp 1
transform 1 0 71392 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input37
timestamp 1
transform -1 0 72680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1
transform -1 0 29992 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input39
timestamp 1
transform 1 0 33764 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1
transform 1 0 35328 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input41
timestamp 1
transform 1 0 36432 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1
transform -1 0 38180 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1
transform -1 0 39192 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input44
timestamp 1
transform -1 0 41768 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  input45
timestamp 1
transform 1 0 27232 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input46
timestamp 1
transform 1 0 28980 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input47
timestamp 1
transform 1 0 30452 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  input48
timestamp 1
transform 1 0 32752 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  input49
timestamp 1
transform 1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input50
timestamp 1
transform 1 0 26864 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output51
timestamp 1
transform -1 0 25760 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output52
timestamp 1
transform -1 0 28244 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 1
transform 1 0 42412 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 1
transform 1 0 43884 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 1
transform 1 0 45172 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 1
transform 1 0 47472 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 1
transform 1 0 47932 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 1
transform 1 0 50048 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 1
transform 1 0 50692 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 1
transform 1 0 52624 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 1
transform 1 0 53452 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 1
transform 1 0 55200 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 1
transform -1 0 29348 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1
transform 1 0 56212 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1
transform 1 0 57592 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1
transform 1 0 57592 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1
transform 1 0 63664 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1
transform 1 0 63664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1
transform 1 0 63664 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1
transform 1 0 64584 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1
transform 1 0 66608 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1
transform 1 0 69368 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1
transform 1 0 69368 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1
transform -1 0 31924 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1
transform 1 0 70656 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1
transform 1 0 71392 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1
transform -1 0 33764 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1
transform 1 0 34132 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1
transform 1 0 35512 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1
transform 1 0 37168 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1
transform 1 0 38180 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1
transform 1 0 39744 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1
transform 1 0 42320 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_0
timestamp 1
transform 1 0 1012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_9
timestamp 1
transform -1 0 74980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_1
timestamp 1
transform 1 0 1012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_10
timestamp 1
transform -1 0 74980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_2
timestamp 1
transform 1 0 1012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_11
timestamp 1
transform -1 0 74980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_3
timestamp 1
transform 1 0 1012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_12
timestamp 1
transform -1 0 74980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_4
timestamp 1
transform 1 0 1012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_13
timestamp 1
transform -1 0 74980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_5
timestamp 1
transform 1 0 1012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_14
timestamp 1
transform -1 0 74980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_6
timestamp 1
transform 1 0 1012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_15
timestamp 1
transform -1 0 74980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_7
timestamp 1
transform 1 0 1012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_16
timestamp 1
transform -1 0 74980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_8
timestamp 1
transform 1 0 1012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_17
timestamp 1
transform -1 0 74980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Left_311
timestamp 1
transform 1 0 65412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Right_164
timestamp 1
transform -1 0 74980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_165
timestamp 1
transform 1 0 65412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_18
timestamp 1
transform -1 0 74980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_166
timestamp 1
transform 1 0 65412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_19
timestamp 1
transform -1 0 74980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_167
timestamp 1
transform 1 0 65412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_20
timestamp 1
transform -1 0 74980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_168
timestamp 1
transform 1 0 65412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_21
timestamp 1
transform -1 0 74980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_169
timestamp 1
transform 1 0 65412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_22
timestamp 1
transform -1 0 74980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_170
timestamp 1
transform 1 0 65412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_23
timestamp 1
transform -1 0 74980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_171
timestamp 1
transform 1 0 65412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_24
timestamp 1
transform -1 0 74980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_172
timestamp 1
transform 1 0 65412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_25
timestamp 1
transform -1 0 74980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_173
timestamp 1
transform 1 0 65412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_26
timestamp 1
transform -1 0 74980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_174
timestamp 1
transform 1 0 65412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_27
timestamp 1
transform -1 0 74980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_175
timestamp 1
transform 1 0 65412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_28
timestamp 1
transform -1 0 74980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_176
timestamp 1
transform 1 0 65412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_29
timestamp 1
transform -1 0 74980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_177
timestamp 1
transform 1 0 65412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_30
timestamp 1
transform -1 0 74980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_178
timestamp 1
transform 1 0 65412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_31
timestamp 1
transform -1 0 74980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_179
timestamp 1
transform 1 0 65412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_32
timestamp 1
transform -1 0 74980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_180
timestamp 1
transform 1 0 65412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_33
timestamp 1
transform -1 0 74980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_181
timestamp 1
transform 1 0 65412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_34
timestamp 1
transform -1 0 74980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_182
timestamp 1
transform 1 0 65412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_35
timestamp 1
transform -1 0 74980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_183
timestamp 1
transform 1 0 65412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_36
timestamp 1
transform -1 0 74980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_184
timestamp 1
transform 1 0 65412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_37
timestamp 1
transform -1 0 74980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_185
timestamp 1
transform 1 0 65412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_38
timestamp 1
transform -1 0 74980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_186
timestamp 1
transform 1 0 65412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_39
timestamp 1
transform -1 0 74980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_187
timestamp 1
transform 1 0 65412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_40
timestamp 1
transform -1 0 74980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_188
timestamp 1
transform 1 0 65412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_41
timestamp 1
transform -1 0 74980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_189
timestamp 1
transform 1 0 65412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_42
timestamp 1
transform -1 0 74980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_190
timestamp 1
transform 1 0 65412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_43
timestamp 1
transform -1 0 74980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_191
timestamp 1
transform 1 0 65412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_44
timestamp 1
transform -1 0 74980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_192
timestamp 1
transform 1 0 65412 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_45
timestamp 1
transform -1 0 74980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_193
timestamp 1
transform 1 0 65412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_46
timestamp 1
transform -1 0 74980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_194
timestamp 1
transform 1 0 65412 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_47
timestamp 1
transform -1 0 74980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_195
timestamp 1
transform 1 0 65412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_48
timestamp 1
transform -1 0 74980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_196
timestamp 1
transform 1 0 65412 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_49
timestamp 1
transform -1 0 74980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_197
timestamp 1
transform 1 0 65412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_50
timestamp 1
transform -1 0 74980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_198
timestamp 1
transform 1 0 65412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_51
timestamp 1
transform -1 0 74980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_199
timestamp 1
transform 1 0 65412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_52
timestamp 1
transform -1 0 74980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_200
timestamp 1
transform 1 0 65412 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_53
timestamp 1
transform -1 0 74980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_201
timestamp 1
transform 1 0 65412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_54
timestamp 1
transform -1 0 74980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_202
timestamp 1
transform 1 0 65412 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_55
timestamp 1
transform -1 0 74980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_203
timestamp 1
transform 1 0 65412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_56
timestamp 1
transform -1 0 74980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_204
timestamp 1
transform 1 0 65412 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_57
timestamp 1
transform -1 0 74980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_205
timestamp 1
transform 1 0 65412 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_58
timestamp 1
transform -1 0 74980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_206
timestamp 1
transform 1 0 65412 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_59
timestamp 1
transform -1 0 74980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_207
timestamp 1
transform 1 0 65412 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_60
timestamp 1
transform -1 0 74980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_208
timestamp 1
transform 1 0 65412 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_61
timestamp 1
transform -1 0 74980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_209
timestamp 1
transform 1 0 65412 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_62
timestamp 1
transform -1 0 74980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_210
timestamp 1
transform 1 0 65412 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_63
timestamp 1
transform -1 0 74980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_211
timestamp 1
transform 1 0 65412 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_64
timestamp 1
transform -1 0 74980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_212
timestamp 1
transform 1 0 65412 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_65
timestamp 1
transform -1 0 74980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_213
timestamp 1
transform 1 0 65412 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_66
timestamp 1
transform -1 0 74980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_214
timestamp 1
transform 1 0 65412 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_67
timestamp 1
transform -1 0 74980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_215
timestamp 1
transform 1 0 65412 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_68
timestamp 1
transform -1 0 74980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_216
timestamp 1
transform 1 0 65412 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_69
timestamp 1
transform -1 0 74980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_217
timestamp 1
transform 1 0 65412 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_70
timestamp 1
transform -1 0 74980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_218
timestamp 1
transform 1 0 65412 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_71
timestamp 1
transform -1 0 74980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_219
timestamp 1
transform 1 0 65412 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_72
timestamp 1
transform -1 0 74980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_220
timestamp 1
transform 1 0 65412 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_73
timestamp 1
transform -1 0 74980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_221
timestamp 1
transform 1 0 65412 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_74
timestamp 1
transform -1 0 74980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_222
timestamp 1
transform 1 0 65412 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_75
timestamp 1
transform -1 0 74980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_223
timestamp 1
transform 1 0 65412 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_76
timestamp 1
transform -1 0 74980 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_224
timestamp 1
transform 1 0 65412 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_77
timestamp 1
transform -1 0 74980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_225
timestamp 1
transform 1 0 65412 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_78
timestamp 1
transform -1 0 74980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_226
timestamp 1
transform 1 0 65412 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_79
timestamp 1
transform -1 0 74980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_227
timestamp 1
transform 1 0 65412 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_80
timestamp 1
transform -1 0 74980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_228
timestamp 1
transform 1 0 65412 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_81
timestamp 1
transform -1 0 74980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_229
timestamp 1
transform 1 0 65412 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_82
timestamp 1
transform -1 0 74980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_230
timestamp 1
transform 1 0 65412 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_83
timestamp 1
transform -1 0 74980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_231
timestamp 1
transform 1 0 65412 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_84
timestamp 1
transform -1 0 74980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_232
timestamp 1
transform 1 0 65412 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_85
timestamp 1
transform -1 0 74980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_233
timestamp 1
transform 1 0 65412 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_86
timestamp 1
transform -1 0 74980 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_234
timestamp 1
transform 1 0 65412 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_87
timestamp 1
transform -1 0 74980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_235
timestamp 1
transform 1 0 65412 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_88
timestamp 1
transform -1 0 74980 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_236
timestamp 1
transform 1 0 65412 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_89
timestamp 1
transform -1 0 74980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_237
timestamp 1
transform 1 0 65412 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_90
timestamp 1
transform -1 0 74980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_238
timestamp 1
transform 1 0 65412 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_91
timestamp 1
transform -1 0 74980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_239
timestamp 1
transform 1 0 65412 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_92
timestamp 1
transform -1 0 74980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_240
timestamp 1
transform 1 0 65412 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_93
timestamp 1
transform -1 0 74980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_241
timestamp 1
transform 1 0 65412 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_94
timestamp 1
transform -1 0 74980 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_242
timestamp 1
transform 1 0 65412 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_95
timestamp 1
transform -1 0 74980 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_243
timestamp 1
transform 1 0 65412 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_96
timestamp 1
transform -1 0 74980 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_244
timestamp 1
transform 1 0 65412 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_97
timestamp 1
transform -1 0 74980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_245
timestamp 1
transform 1 0 65412 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_98
timestamp 1
transform -1 0 74980 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_246
timestamp 1
transform 1 0 65412 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_99
timestamp 1
transform -1 0 74980 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_247
timestamp 1
transform 1 0 65412 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_100
timestamp 1
transform -1 0 74980 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_248
timestamp 1
transform 1 0 65412 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_101
timestamp 1
transform -1 0 74980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_249
timestamp 1
transform 1 0 65412 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_102
timestamp 1
transform -1 0 74980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_250
timestamp 1
transform 1 0 65412 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_103
timestamp 1
transform -1 0 74980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_251
timestamp 1
transform 1 0 65412 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_104
timestamp 1
transform -1 0 74980 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_252
timestamp 1
transform 1 0 65412 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_105
timestamp 1
transform -1 0 74980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_253
timestamp 1
transform 1 0 65412 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_106
timestamp 1
transform -1 0 74980 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_254
timestamp 1
transform 1 0 65412 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_107
timestamp 1
transform -1 0 74980 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_255
timestamp 1
transform 1 0 65412 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_108
timestamp 1
transform -1 0 74980 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_256
timestamp 1
transform 1 0 65412 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_109
timestamp 1
transform -1 0 74980 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_257
timestamp 1
transform 1 0 65412 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_110
timestamp 1
transform -1 0 74980 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_258
timestamp 1
transform 1 0 65412 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_111
timestamp 1
transform -1 0 74980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_259
timestamp 1
transform 1 0 65412 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_112
timestamp 1
transform -1 0 74980 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_260
timestamp 1
transform 1 0 65412 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_113
timestamp 1
transform -1 0 74980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Left_261
timestamp 1
transform 1 0 65412 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_2_Right_114
timestamp 1
transform -1 0 74980 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Left_262
timestamp 1
transform 1 0 65412 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_2_Right_115
timestamp 1
transform -1 0 74980 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Left_263
timestamp 1
transform 1 0 65412 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_2_Right_116
timestamp 1
transform -1 0 74980 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Left_264
timestamp 1
transform 1 0 65412 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_2_Right_117
timestamp 1
transform -1 0 74980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Left_265
timestamp 1
transform 1 0 65412 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_2_Right_118
timestamp 1
transform -1 0 74980 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Left_266
timestamp 1
transform 1 0 65412 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_2_Right_119
timestamp 1
transform -1 0 74980 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Left_267
timestamp 1
transform 1 0 65412 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_2_Right_120
timestamp 1
transform -1 0 74980 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Left_268
timestamp 1
transform 1 0 65412 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_2_Right_121
timestamp 1
transform -1 0 74980 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Left_269
timestamp 1
transform 1 0 65412 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_2_Right_122
timestamp 1
transform -1 0 74980 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Left_270
timestamp 1
transform 1 0 65412 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_2_Right_123
timestamp 1
transform -1 0 74980 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Left_271
timestamp 1
transform 1 0 65412 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_2_Right_124
timestamp 1
transform -1 0 74980 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Left_272
timestamp 1
transform 1 0 65412 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_2_Right_125
timestamp 1
transform -1 0 74980 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Left_273
timestamp 1
transform 1 0 65412 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_2_Right_126
timestamp 1
transform -1 0 74980 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Left_274
timestamp 1
transform 1 0 65412 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_2_Right_127
timestamp 1
transform -1 0 74980 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Left_275
timestamp 1
transform 1 0 65412 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_2_Right_128
timestamp 1
transform -1 0 74980 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Left_276
timestamp 1
transform 1 0 65412 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_2_Right_129
timestamp 1
transform -1 0 74980 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Left_277
timestamp 1
transform 1 0 65412 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_2_Right_130
timestamp 1
transform -1 0 74980 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Left_278
timestamp 1
transform 1 0 65412 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_2_Right_131
timestamp 1
transform -1 0 74980 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Left_279
timestamp 1
transform 1 0 65412 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_2_Right_132
timestamp 1
transform -1 0 74980 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Left_280
timestamp 1
transform 1 0 65412 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_2_Right_133
timestamp 1
transform -1 0 74980 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Left_281
timestamp 1
transform 1 0 65412 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_2_Right_134
timestamp 1
transform -1 0 74980 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Left_282
timestamp 1
transform 1 0 65412 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_2_Right_135
timestamp 1
transform -1 0 74980 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Left_283
timestamp 1
transform 1 0 65412 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_2_Right_136
timestamp 1
transform -1 0 74980 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Left_284
timestamp 1
transform 1 0 65412 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_2_Right_137
timestamp 1
transform -1 0 74980 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Left_285
timestamp 1
transform 1 0 65412 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_2_Right_138
timestamp 1
transform -1 0 74980 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Left_286
timestamp 1
transform 1 0 65412 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_2_Right_139
timestamp 1
transform -1 0 74980 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Left_287
timestamp 1
transform 1 0 65412 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_2_Right_140
timestamp 1
transform -1 0 74980 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Left_288
timestamp 1
transform 1 0 65412 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_2_Right_141
timestamp 1
transform -1 0 74980 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Left_289
timestamp 1
transform 1 0 65412 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_2_Right_142
timestamp 1
transform -1 0 74980 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Left_290
timestamp 1
transform 1 0 65412 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_2_Right_143
timestamp 1
transform -1 0 74980 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Left_291
timestamp 1
transform 1 0 65412 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_2_Right_144
timestamp 1
transform -1 0 74980 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Left_292
timestamp 1
transform 1 0 65412 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_2_Right_145
timestamp 1
transform -1 0 74980 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Left_293
timestamp 1
transform 1 0 65412 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_2_Right_146
timestamp 1
transform -1 0 74980 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Left_294
timestamp 1
transform 1 0 65412 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_2_Right_147
timestamp 1
transform -1 0 74980 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Left_295
timestamp 1
transform 1 0 65412 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_2_Right_148
timestamp 1
transform -1 0 74980 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Left_296
timestamp 1
transform 1 0 65412 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_2_Right_149
timestamp 1
transform -1 0 74980 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Left_297
timestamp 1
transform 1 0 65412 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_2_Right_150
timestamp 1
transform -1 0 74980 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Left_298
timestamp 1
transform 1 0 65412 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_2_Right_151
timestamp 1
transform -1 0 74980 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Left_299
timestamp 1
transform 1 0 65412 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_2_Right_152
timestamp 1
transform -1 0 74980 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Left_300
timestamp 1
transform 1 0 65412 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_2_Right_153
timestamp 1
transform -1 0 74980 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Left_301
timestamp 1
transform 1 0 65412 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_2_Right_154
timestamp 1
transform -1 0 74980 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Left_302
timestamp 1
transform 1 0 65412 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_2_Right_155
timestamp 1
transform -1 0 74980 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Left_303
timestamp 1
transform 1 0 65412 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_2_Right_156
timestamp 1
transform -1 0 74980 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Left_304
timestamp 1
transform 1 0 65412 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_2_Right_157
timestamp 1
transform -1 0 74980 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Left_305
timestamp 1
transform 1 0 65412 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_2_Right_158
timestamp 1
transform -1 0 74980 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Left_306
timestamp 1
transform 1 0 65412 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_2_Right_159
timestamp 1
transform -1 0 74980 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Left_307
timestamp 1
transform 1 0 65412 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_2_Right_160
timestamp 1
transform -1 0 74980 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Left_308
timestamp 1
transform 1 0 65412 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_2_Right_161
timestamp 1
transform -1 0 74980 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Left_309
timestamp 1
transform 1 0 65412 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_2_Right_162
timestamp 1
transform -1 0 74980 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Left_310
timestamp 1
transform 1 0 65412 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_2_Right_163
timestamp 1
transform -1 0 74980 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_312
timestamp 1
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_313
timestamp 1
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_314
timestamp 1
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_315
timestamp 1
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_316
timestamp 1
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_317
timestamp 1
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_318
timestamp 1
transform 1 0 19044 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_319
timestamp 1
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_320
timestamp 1
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_321
timestamp 1
transform 1 0 26772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_322
timestamp 1
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_323
timestamp 1
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_324
timestamp 1
transform 1 0 34500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_325
timestamp 1
transform 1 0 37076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_326
timestamp 1
transform 1 0 39652 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_327
timestamp 1
transform 1 0 42228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_328
timestamp 1
transform 1 0 44804 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_329
timestamp 1
transform 1 0 47380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_330
timestamp 1
transform 1 0 49956 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_331
timestamp 1
transform 1 0 52532 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_332
timestamp 1
transform 1 0 55108 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_333
timestamp 1
transform 1 0 57684 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_334
timestamp 1
transform 1 0 60260 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_335
timestamp 1
transform 1 0 62836 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_336
timestamp 1
transform 1 0 65412 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_337
timestamp 1
transform 1 0 67988 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_338
timestamp 1
transform 1 0 70564 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_339
timestamp 1
transform 1 0 73140 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_340
timestamp 1
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_341
timestamp 1
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_342
timestamp 1
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_343
timestamp 1
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_344
timestamp 1
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_345
timestamp 1
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_346
timestamp 1
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_347
timestamp 1
transform 1 0 42228 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_348
timestamp 1
transform 1 0 47380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_349
timestamp 1
transform 1 0 52532 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_350
timestamp 1
transform 1 0 57684 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_351
timestamp 1
transform 1 0 62836 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_352
timestamp 1
transform 1 0 67988 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_353
timestamp 1
transform 1 0 73140 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_354
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_355
timestamp 1
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_356
timestamp 1
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_357
timestamp 1
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_358
timestamp 1
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_359
timestamp 1
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_360
timestamp 1
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_361
timestamp 1
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_362
timestamp 1
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_363
timestamp 1
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_364
timestamp 1
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_365
timestamp 1
transform 1 0 60260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_366
timestamp 1
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_367
timestamp 1
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_368
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_369
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_370
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_371
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_372
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_373
timestamp 1
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_374
timestamp 1
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_375
timestamp 1
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_376
timestamp 1
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_377
timestamp 1
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_378
timestamp 1
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_379
timestamp 1
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_380
timestamp 1
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_381
timestamp 1
transform 1 0 73140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_382
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_383
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_384
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_385
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_386
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_387
timestamp 1
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_388
timestamp 1
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_389
timestamp 1
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_390
timestamp 1
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_391
timestamp 1
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_392
timestamp 1
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_393
timestamp 1
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_394
timestamp 1
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_395
timestamp 1
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_396
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_397
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_398
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_399
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_400
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_401
timestamp 1
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_402
timestamp 1
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_403
timestamp 1
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_404
timestamp 1
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_405
timestamp 1
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_406
timestamp 1
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_407
timestamp 1
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_408
timestamp 1
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_409
timestamp 1
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_410
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_411
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_412
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_413
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_414
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_415
timestamp 1
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_416
timestamp 1
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_417
timestamp 1
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_418
timestamp 1
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_419
timestamp 1
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_420
timestamp 1
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_421
timestamp 1
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_422
timestamp 1
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_423
timestamp 1
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_424
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_425
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_426
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_427
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_428
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_429
timestamp 1
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_430
timestamp 1
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_431
timestamp 1
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_432
timestamp 1
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_433
timestamp 1
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_434
timestamp 1
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_435
timestamp 1
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_436
timestamp 1
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_437
timestamp 1
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_438
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_439
timestamp 1
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_440
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_441
timestamp 1
transform 1 0 11316 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_442
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_443
timestamp 1
transform 1 0 16468 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_444
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_445
timestamp 1
transform 1 0 21620 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_446
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_447
timestamp 1
transform 1 0 26772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_448
timestamp 1
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_449
timestamp 1
transform 1 0 31924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_450
timestamp 1
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_451
timestamp 1
transform 1 0 37076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_452
timestamp 1
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_453
timestamp 1
transform 1 0 42228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_454
timestamp 1
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_455
timestamp 1
transform 1 0 47380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_456
timestamp 1
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_457
timestamp 1
transform 1 0 52532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_458
timestamp 1
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_459
timestamp 1
transform 1 0 57684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_460
timestamp 1
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_461
timestamp 1
transform 1 0 62836 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_462
timestamp 1
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_463
timestamp 1
transform 1 0 67988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_464
timestamp 1
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_465
timestamp 1
transform 1 0 73140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_2_687
timestamp 1
transform 1 0 70564 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_466
timestamp 1
transform 1 0 67988 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_467
timestamp 1
transform 1 0 73140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_468
timestamp 1
transform 1 0 70564 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_469
timestamp 1
transform 1 0 67988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_470
timestamp 1
transform 1 0 73140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_471
timestamp 1
transform 1 0 70564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_472
timestamp 1
transform 1 0 67988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_2_473
timestamp 1
transform 1 0 73140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_2_474
timestamp 1
transform 1 0 70564 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_475
timestamp 1
transform 1 0 67988 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_2_476
timestamp 1
transform 1 0 73140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_2_477
timestamp 1
transform 1 0 70564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_478
timestamp 1
transform 1 0 67988 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_2_479
timestamp 1
transform 1 0 73140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_2_480
timestamp 1
transform 1 0 70564 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_481
timestamp 1
transform 1 0 67988 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_2_482
timestamp 1
transform 1 0 73140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_2_483
timestamp 1
transform 1 0 70564 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_484
timestamp 1
transform 1 0 67988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_2_485
timestamp 1
transform 1 0 73140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_2_486
timestamp 1
transform 1 0 70564 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_487
timestamp 1
transform 1 0 67988 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_2_488
timestamp 1
transform 1 0 73140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_2_489
timestamp 1
transform 1 0 70564 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_490
timestamp 1
transform 1 0 67988 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_2_491
timestamp 1
transform 1 0 73140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_2_492
timestamp 1
transform 1 0 70564 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_493
timestamp 1
transform 1 0 67988 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_2_494
timestamp 1
transform 1 0 73140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_2_495
timestamp 1
transform 1 0 70564 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_496
timestamp 1
transform 1 0 67988 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_2_497
timestamp 1
transform 1 0 73140 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_2_498
timestamp 1
transform 1 0 70564 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_499
timestamp 1
transform 1 0 67988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_2_500
timestamp 1
transform 1 0 73140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_2_501
timestamp 1
transform 1 0 70564 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_502
timestamp 1
transform 1 0 67988 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_2_503
timestamp 1
transform 1 0 73140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_2_504
timestamp 1
transform 1 0 70564 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_505
timestamp 1
transform 1 0 67988 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_2_506
timestamp 1
transform 1 0 73140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_2_507
timestamp 1
transform 1 0 70564 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_508
timestamp 1
transform 1 0 67988 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_2_509
timestamp 1
transform 1 0 73140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_2_510
timestamp 1
transform 1 0 70564 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_511
timestamp 1
transform 1 0 67988 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_2_512
timestamp 1
transform 1 0 73140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_2_513
timestamp 1
transform 1 0 70564 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_514
timestamp 1
transform 1 0 67988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_2_515
timestamp 1
transform 1 0 73140 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_2_516
timestamp 1
transform 1 0 70564 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_517
timestamp 1
transform 1 0 67988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_2_518
timestamp 1
transform 1 0 73140 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_2_519
timestamp 1
transform 1 0 70564 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_520
timestamp 1
transform 1 0 67988 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_2_521
timestamp 1
transform 1 0 73140 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_2_522
timestamp 1
transform 1 0 70564 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_523
timestamp 1
transform 1 0 67988 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_2_524
timestamp 1
transform 1 0 73140 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_2_525
timestamp 1
transform 1 0 70564 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_526
timestamp 1
transform 1 0 67988 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_2_527
timestamp 1
transform 1 0 73140 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_2_528
timestamp 1
transform 1 0 70564 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_529
timestamp 1
transform 1 0 67988 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_2_530
timestamp 1
transform 1 0 73140 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_2_531
timestamp 1
transform 1 0 70564 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_532
timestamp 1
transform 1 0 67988 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_2_533
timestamp 1
transform 1 0 73140 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_2_534
timestamp 1
transform 1 0 70564 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_535
timestamp 1
transform 1 0 67988 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_2_536
timestamp 1
transform 1 0 73140 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_2_537
timestamp 1
transform 1 0 70564 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_538
timestamp 1
transform 1 0 67988 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_2_539
timestamp 1
transform 1 0 73140 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_2_540
timestamp 1
transform 1 0 70564 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_541
timestamp 1
transform 1 0 67988 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_2_542
timestamp 1
transform 1 0 73140 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_2_543
timestamp 1
transform 1 0 70564 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_544
timestamp 1
transform 1 0 67988 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_2_545
timestamp 1
transform 1 0 73140 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_2_546
timestamp 1
transform 1 0 70564 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_547
timestamp 1
transform 1 0 67988 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_2_548
timestamp 1
transform 1 0 73140 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_2_549
timestamp 1
transform 1 0 70564 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_550
timestamp 1
transform 1 0 67988 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_2_551
timestamp 1
transform 1 0 73140 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_2_552
timestamp 1
transform 1 0 70564 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_553
timestamp 1
transform 1 0 67988 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_2_554
timestamp 1
transform 1 0 73140 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_2_555
timestamp 1
transform 1 0 70564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_556
timestamp 1
transform 1 0 67988 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_2_557
timestamp 1
transform 1 0 73140 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_2_558
timestamp 1
transform 1 0 70564 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_559
timestamp 1
transform 1 0 67988 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_2_560
timestamp 1
transform 1 0 73140 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_2_561
timestamp 1
transform 1 0 70564 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_562
timestamp 1
transform 1 0 67988 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_2_563
timestamp 1
transform 1 0 73140 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_2_564
timestamp 1
transform 1 0 70564 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_565
timestamp 1
transform 1 0 67988 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_2_566
timestamp 1
transform 1 0 73140 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_2_567
timestamp 1
transform 1 0 70564 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_568
timestamp 1
transform 1 0 67988 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_2_569
timestamp 1
transform 1 0 73140 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_2_570
timestamp 1
transform 1 0 70564 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_571
timestamp 1
transform 1 0 67988 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_2_572
timestamp 1
transform 1 0 73140 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_2_573
timestamp 1
transform 1 0 70564 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_574
timestamp 1
transform 1 0 67988 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_2_575
timestamp 1
transform 1 0 73140 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_2_576
timestamp 1
transform 1 0 70564 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_577
timestamp 1
transform 1 0 67988 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_2_578
timestamp 1
transform 1 0 73140 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_2_579
timestamp 1
transform 1 0 70564 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_580
timestamp 1
transform 1 0 67988 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_2_581
timestamp 1
transform 1 0 73140 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_2_582
timestamp 1
transform 1 0 70564 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_583
timestamp 1
transform 1 0 67988 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_2_584
timestamp 1
transform 1 0 73140 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_2_585
timestamp 1
transform 1 0 70564 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_586
timestamp 1
transform 1 0 67988 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_2_587
timestamp 1
transform 1 0 73140 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_2_588
timestamp 1
transform 1 0 70564 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_589
timestamp 1
transform 1 0 67988 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_2_590
timestamp 1
transform 1 0 73140 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_2_591
timestamp 1
transform 1 0 70564 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_592
timestamp 1
transform 1 0 67988 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_2_593
timestamp 1
transform 1 0 73140 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_2_594
timestamp 1
transform 1 0 70564 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_595
timestamp 1
transform 1 0 67988 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_2_596
timestamp 1
transform 1 0 73140 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_2_597
timestamp 1
transform 1 0 70564 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_598
timestamp 1
transform 1 0 67988 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_2_599
timestamp 1
transform 1 0 73140 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_2_600
timestamp 1
transform 1 0 70564 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_601
timestamp 1
transform 1 0 67988 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_2_602
timestamp 1
transform 1 0 73140 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_2_603
timestamp 1
transform 1 0 70564 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_604
timestamp 1
transform 1 0 67988 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_2_605
timestamp 1
transform 1 0 73140 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_2_606
timestamp 1
transform 1 0 70564 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_607
timestamp 1
transform 1 0 67988 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_2_608
timestamp 1
transform 1 0 73140 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_2_609
timestamp 1
transform 1 0 70564 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_610
timestamp 1
transform 1 0 67988 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_2_611
timestamp 1
transform 1 0 73140 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_2_612
timestamp 1
transform 1 0 70564 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_613
timestamp 1
transform 1 0 67988 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_2_614
timestamp 1
transform 1 0 73140 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_2_615
timestamp 1
transform 1 0 70564 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_616
timestamp 1
transform 1 0 67988 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_2_617
timestamp 1
transform 1 0 73140 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_2_618
timestamp 1
transform 1 0 70564 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_619
timestamp 1
transform 1 0 67988 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_2_620
timestamp 1
transform 1 0 73140 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_2_621
timestamp 1
transform 1 0 70564 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_622
timestamp 1
transform 1 0 67988 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_2_623
timestamp 1
transform 1 0 73140 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_2_624
timestamp 1
transform 1 0 70564 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_625
timestamp 1
transform 1 0 67988 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_2_626
timestamp 1
transform 1 0 73140 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2_627
timestamp 1
transform 1 0 70564 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_628
timestamp 1
transform 1 0 67988 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2_629
timestamp 1
transform 1 0 73140 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2_630
timestamp 1
transform 1 0 70564 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_631
timestamp 1
transform 1 0 67988 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2_632
timestamp 1
transform 1 0 73140 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2_633
timestamp 1
transform 1 0 70564 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_634
timestamp 1
transform 1 0 67988 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2_635
timestamp 1
transform 1 0 73140 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2_636
timestamp 1
transform 1 0 70564 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_637
timestamp 1
transform 1 0 67988 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2_638
timestamp 1
transform 1 0 73140 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2_639
timestamp 1
transform 1 0 70564 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_640
timestamp 1
transform 1 0 67988 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2_641
timestamp 1
transform 1 0 73140 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2_642
timestamp 1
transform 1 0 70564 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_643
timestamp 1
transform 1 0 67988 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2_644
timestamp 1
transform 1 0 73140 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2_645
timestamp 1
transform 1 0 70564 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_646
timestamp 1
transform 1 0 67988 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2_647
timestamp 1
transform 1 0 73140 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2_648
timestamp 1
transform 1 0 70564 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_649
timestamp 1
transform 1 0 67988 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2_650
timestamp 1
transform 1 0 73140 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2_651
timestamp 1
transform 1 0 70564 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_652
timestamp 1
transform 1 0 67988 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2_653
timestamp 1
transform 1 0 73140 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2_654
timestamp 1
transform 1 0 70564 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_655
timestamp 1
transform 1 0 67988 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2_656
timestamp 1
transform 1 0 73140 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2_657
timestamp 1
transform 1 0 70564 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_658
timestamp 1
transform 1 0 67988 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2_659
timestamp 1
transform 1 0 73140 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_2_660
timestamp 1
transform 1 0 70564 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_661
timestamp 1
transform 1 0 67988 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_2_662
timestamp 1
transform 1 0 73140 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_2_663
timestamp 1
transform 1 0 70564 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_664
timestamp 1
transform 1 0 67988 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_2_665
timestamp 1
transform 1 0 73140 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_2_666
timestamp 1
transform 1 0 70564 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_667
timestamp 1
transform 1 0 67988 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_2_668
timestamp 1
transform 1 0 73140 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_2_669
timestamp 1
transform 1 0 70564 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_670
timestamp 1
transform 1 0 67988 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_2_671
timestamp 1
transform 1 0 73140 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_2_672
timestamp 1
transform 1 0 70564 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_673
timestamp 1
transform 1 0 67988 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_2_674
timestamp 1
transform 1 0 73140 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_2_675
timestamp 1
transform 1 0 70564 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_676
timestamp 1
transform 1 0 67988 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_2_677
timestamp 1
transform 1 0 73140 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_2_678
timestamp 1
transform 1 0 70564 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_679
timestamp 1
transform 1 0 67988 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_2_680
timestamp 1
transform 1 0 73140 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_2_681
timestamp 1
transform 1 0 70564 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_682
timestamp 1
transform 1 0 67988 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_2_683
timestamp 1
transform 1 0 73140 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_684
timestamp 1
transform 1 0 67988 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_685
timestamp 1
transform 1 0 70564 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_2_686
timestamp 1
transform 1 0 73140 0 -1 85952
box -38 -48 130 592
<< labels >>
flabel metal2 s 4188 1040 4540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 14188 1040 14540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 24188 1040 24540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 34188 1040 34540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 44188 1040 44540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 54188 1040 54540 5944 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 64188 1040 64540 5972 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 74188 1040 74540 86000 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 4264 75028 4616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 14264 75028 14616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 24264 75028 24616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 34264 75028 34616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 44264 75028 44616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 54264 75028 54616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 64264 75028 64616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 74264 75028 74616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 964 84264 75028 84616 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4702 0 5322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4702 0 5322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4702 86940 5322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10702 0 11322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10702 0 11322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10702 86940 11322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16702 0 17322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16702 0 17322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16702 86940 17322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 22702 0 23322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 22702 0 23322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 22702 86940 23322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 28702 0 29322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 28702 0 29322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 28702 86940 29322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 34702 0 35322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 34702 0 35322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 34702 86940 35322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 40702 0 41322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 40702 0 41322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 40702 86940 41322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 46702 0 47322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 46702 0 47322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 46702 86940 47322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 52702 0 53322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 52702 0 53322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 52702 86940 53322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 58702 0 59322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 58702 0 59322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 58702 86940 59322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 64702 0 65322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 64702 0 65322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 64702 86940 65322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 70702 0 71322 87000 0 FreeSans 3840 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 70702 0 71322 60 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 70702 86940 71322 87000 0 FreeSans 480 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 1836 1040 2188 5944 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 11836 1040 12188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 21836 1040 22188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 31836 1040 32188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 41836 1040 42188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 51836 1040 52188 5944 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 61836 1040 62188 5972 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 71836 1040 72188 86000 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 1912 75028 2264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 11912 75028 12264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 21912 75028 22264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 31912 75028 32264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 41912 75028 42264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 51912 75028 52264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 61912 75028 62264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 71912 75028 72264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 964 81912 75028 82264 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 1702 0 2322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 1702 0 2322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 1702 86940 2322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7702 0 8322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7702 0 8322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7702 86940 8322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13702 0 14322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13702 0 14322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13702 86940 14322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19702 0 20322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19702 0 20322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19702 86940 20322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 25702 0 26322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 25702 0 26322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 25702 86940 26322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 31702 0 32322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 31702 0 32322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 31702 86940 32322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 37702 0 38322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 37702 0 38322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 37702 86940 38322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 43702 0 44322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 43702 0 44322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 43702 86940 44322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 49702 0 50322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 49702 0 50322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 49702 86940 50322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 55702 0 56322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 55702 0 56322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 55702 86940 56322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 61702 0 62322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 61702 0 62322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 61702 86940 62322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 67702 0 68322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 67702 0 68322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 67702 86940 68322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 73702 0 74322 87000 0 FreeSans 3840 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 73702 0 74322 60 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 73702 86940 74322 87000 0 FreeSans 480 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 wb_clk_i
port 2 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 wb_rst_i
port 3 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 4 nsew signal output
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 5 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 6 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 7 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 8 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 9 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 10 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 11 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 12 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 13 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 14 nsew signal input
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 15 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 16 nsew signal input
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 17 nsew signal input
flabel metal2 s 56598 0 56654 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 18 nsew signal input
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 19 nsew signal input
flabel metal2 s 59358 0 59414 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 20 nsew signal input
flabel metal2 s 60738 0 60794 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 21 nsew signal input
flabel metal2 s 62118 0 62174 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 22 nsew signal input
flabel metal2 s 63498 0 63554 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 23 nsew signal input
flabel metal2 s 64878 0 64934 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 24 nsew signal input
flabel metal2 s 66258 0 66314 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 25 nsew signal input
flabel metal2 s 67638 0 67694 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 26 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 27 nsew signal input
flabel metal2 s 69018 0 69074 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 28 nsew signal input
flabel metal2 s 70398 0 70454 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 29 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 30 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 31 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 32 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 33 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 34 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 35 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 36 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 37 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 38 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 39 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 40 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 41 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 42 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 43 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 44 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 45 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 46 nsew signal input
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 47 nsew signal input
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 48 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 49 nsew signal input
flabel metal2 s 55678 0 55734 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 50 nsew signal input
flabel metal2 s 57058 0 57114 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 51 nsew signal input
flabel metal2 s 58438 0 58494 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 52 nsew signal input
flabel metal2 s 59818 0 59874 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 53 nsew signal input
flabel metal2 s 61198 0 61254 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 54 nsew signal input
flabel metal2 s 62578 0 62634 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 55 nsew signal input
flabel metal2 s 63958 0 64014 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 56 nsew signal input
flabel metal2 s 65338 0 65394 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 57 nsew signal input
flabel metal2 s 66718 0 66774 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 58 nsew signal input
flabel metal2 s 68098 0 68154 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 59 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 60 nsew signal input
flabel metal2 s 69478 0 69534 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 61 nsew signal input
flabel metal2 s 70858 0 70914 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 62 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 63 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 64 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 65 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 66 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 67 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 68 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 69 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 70 nsew signal output
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 71 nsew signal output
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 72 nsew signal output
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 73 nsew signal output
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 74 nsew signal output
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 75 nsew signal output
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 76 nsew signal output
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 77 nsew signal output
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 78 nsew signal output
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 79 nsew signal output
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 80 nsew signal output
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 81 nsew signal output
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 82 nsew signal output
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 83 nsew signal output
flabel metal2 s 58898 0 58954 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 84 nsew signal output
flabel metal2 s 60278 0 60334 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 85 nsew signal output
flabel metal2 s 61658 0 61714 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 86 nsew signal output
flabel metal2 s 63038 0 63094 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 87 nsew signal output
flabel metal2 s 64418 0 64474 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 88 nsew signal output
flabel metal2 s 65798 0 65854 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 89 nsew signal output
flabel metal2 s 67178 0 67234 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 90 nsew signal output
flabel metal2 s 68558 0 68614 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 91 nsew signal output
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 92 nsew signal output
flabel metal2 s 69938 0 69994 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 93 nsew signal output
flabel metal2 s 71318 0 71374 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 94 nsew signal output
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 95 nsew signal output
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 96 nsew signal output
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 97 nsew signal output
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 98 nsew signal output
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 99 nsew signal output
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 100 nsew signal output
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 101 nsew signal output
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 102 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 103 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 104 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 105 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 106 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 wbs_we_i
port 107 nsew signal input
rlabel via2 62728 84560 62728 84560 0 VGND
rlabel via2 62526 82208 62526 82208 0 VPWR
rlabel metal2 28474 2176 28474 2176 0 _00_
rlabel metal2 47334 5712 47334 5712 0 clknet_0_wb_clk_i
rlabel metal1 35742 3060 35742 3060 0 clknet_1_0__leaf_wb_clk_i
rlabel metal1 63342 53280 63342 53280 0 clknet_1_1__leaf_wb_clk_i
rlabel metal1 63342 43283 63342 43283 0 i_ram_wb_controller.DO\[0\]
rlabel metal1 63342 21421 63342 21421 0 i_ram_wb_controller.DO\[10\]
rlabel metal1 43930 2958 43930 2958 0 i_ram_wb_controller.DO\[11\]
rlabel metal1 63342 17031 63342 17031 0 i_ram_wb_controller.DO\[12\]
rlabel metal1 63342 14853 63342 14853 0 i_ram_wb_controller.DO\[13\]
rlabel metal1 63342 12675 63342 12675 0 i_ram_wb_controller.DO\[14\]
rlabel metal1 53958 4488 53958 4488 0 i_ram_wb_controller.DO\[15\]
rlabel metal1 63250 50288 63250 50288 0 i_ram_wb_controller.DO\[16\]
rlabel metal1 63250 52466 63250 52466 0 i_ram_wb_controller.DO\[17\]
rlabel metal1 63250 54644 63250 54644 0 i_ram_wb_controller.DO\[18\]
rlabel metal1 63342 56754 63342 56754 0 i_ram_wb_controller.DO\[19\]
rlabel metal1 63342 41023 63342 41023 0 i_ram_wb_controller.DO\[1\]
rlabel metal1 63342 58864 63342 58864 0 i_ram_wb_controller.DO\[20\]
rlabel via1 55074 4046 55074 4046 0 i_ram_wb_controller.DO\[21\]
rlabel via1 56546 4046 56546 4046 0 i_ram_wb_controller.DO\[22\]
rlabel via1 58294 4046 58294 4046 0 i_ram_wb_controller.DO\[23\]
rlabel metal1 64400 12002 64400 12002 0 i_ram_wb_controller.DO\[24\]
rlabel metal1 63342 69754 63342 69754 0 i_ram_wb_controller.DO\[25\]
rlabel metal1 63342 72116 63342 72116 0 i_ram_wb_controller.DO\[26\]
rlabel metal1 63342 74110 63342 74110 0 i_ram_wb_controller.DO\[27\]
rlabel metal1 63986 44710 63986 44710 0 i_ram_wb_controller.DO\[28\]
rlabel metal1 63342 78534 63342 78534 0 i_ram_wb_controller.DO\[29\]
rlabel metal1 63342 38811 63342 38811 0 i_ram_wb_controller.DO\[2\]
rlabel metal1 63342 80712 63342 80712 0 i_ram_wb_controller.DO\[30\]
rlabel metal1 63441 83004 63441 83004 0 i_ram_wb_controller.DO\[31\]
rlabel metal1 63342 36633 63342 36633 0 i_ram_wb_controller.DO\[3\]
rlabel metal1 63342 34571 63342 34571 0 i_ram_wb_controller.DO\[4\]
rlabel metal1 63342 32393 63342 32393 0 i_ram_wb_controller.DO\[5\]
rlabel via1 34098 3434 34098 3434 0 i_ram_wb_controller.DO\[6\]
rlabel metal2 32982 5882 32982 5882 0 i_ram_wb_controller.DO\[7\]
rlabel metal2 32614 3553 32614 3553 0 i_ram_wb_controller.DO\[8\]
rlabel via1 31706 4046 31706 4046 0 i_ram_wb_controller.DO\[9\]
rlabel metal1 63986 48790 63986 48790 0 i_ram_wb_controller.EN
rlabel metal1 63342 48105 63342 48105 0 i_ram_wb_controller.R_WB
rlabel metal2 27646 1768 27646 1768 0 net1
rlabel metal2 38870 3196 38870 3196 0 net10
rlabel metal2 57362 6443 57362 6443 0 net100
rlabel metal1 29486 3468 29486 3468 0 net101
rlabel metal1 63625 38658 63625 38658 0 net102
rlabel metal1 42274 3026 42274 3026 0 net103
rlabel metal1 63441 21218 63441 21218 0 net104
rlabel metal1 67344 1938 67344 1938 0 net105
rlabel metal1 63342 74556 63342 74556 0 net106
rlabel metal2 26726 2550 26726 2550 0 net107
rlabel metal1 63342 40829 63342 40829 0 net108
rlabel metal1 67942 2822 67942 2822 0 net109
rlabel metal2 60122 2142 60122 2142 0 net11
rlabel metal1 63441 76716 63441 76716 0 net110
rlabel metal2 41630 3026 41630 3026 0 net111
rlabel metal2 53314 5984 53314 5984 0 net112
rlabel metal1 25484 2074 25484 2074 0 net113
rlabel metal1 63342 42905 63342 42905 0 net114
rlabel metal1 48392 1326 48392 1326 0 net115
rlabel metal2 56626 5950 56626 5950 0 net116
rlabel metal2 70886 2108 70886 2108 0 net117
rlabel metal1 63342 78796 63342 78796 0 net118
rlabel metal2 47058 2108 47058 2108 0 net119
rlabel metal1 24426 2040 24426 2040 0 net12
rlabel metal1 58282 5848 58282 5848 0 net120
rlabel metal1 39146 1938 39146 1938 0 net121
rlabel metal1 52256 5882 52256 5882 0 net122
rlabel metal1 71392 2414 71392 2414 0 net123
rlabel metal1 63342 81008 63342 81008 0 net124
rlabel metal1 45816 2414 45816 2414 0 net125
rlabel metal1 63342 16735 63342 16735 0 net126
rlabel metal1 72956 1258 72956 1258 0 net127
rlabel metal1 63342 83186 63342 83186 0 net128
rlabel metal2 38410 3230 38410 3230 0 net129
rlabel metal2 36478 5168 36478 5168 0 net13
rlabel metal1 54878 5032 54878 5032 0 net130
rlabel metal1 36432 2074 36432 2074 0 net131
rlabel metal2 51474 6256 51474 6256 0 net132
rlabel metal1 45120 3026 45120 3026 0 net133
rlabel metal1 57730 5780 57730 5780 0 net134
rlabel metal1 34040 2278 34040 2278 0 net135
rlabel metal1 63342 31947 63342 31947 0 net136
rlabel metal1 54326 2346 54326 2346 0 net137
rlabel metal1 63342 54838 63342 54838 0 net138
rlabel metal1 44620 2618 44620 2618 0 net139
rlabel metal2 52762 4522 52762 4522 0 net14
rlabel metal1 63342 44309 63342 44309 0 net140
rlabel metal1 52394 2346 52394 2346 0 net141
rlabel metal1 63342 52694 63342 52694 0 net142
rlabel metal2 55798 2108 55798 2108 0 net143
rlabel metal1 63342 57016 63342 57016 0 net144
rlabel metal1 33764 2618 33764 2618 0 net145
rlabel metal1 63342 34125 63342 34125 0 net146
rlabel metal2 50554 1564 50554 1564 0 net147
rlabel metal1 63342 50482 63342 50482 0 net148
rlabel metal1 56994 2346 56994 2346 0 net149
rlabel metal2 51198 4403 51198 4403 0 net15
rlabel metal1 63342 59194 63342 59194 0 net150
rlabel metal1 41676 3026 41676 3026 0 net151
rlabel metal1 63618 37842 63618 37842 0 net152
rlabel metal1 58742 3026 58742 3026 0 net153
rlabel metal1 64492 55250 64492 55250 0 net154
rlabel metal1 59570 2074 59570 2074 0 net155
rlabel metal2 65228 39916 65228 39916 0 net156
rlabel metal1 61226 2346 61226 2346 0 net157
rlabel metal2 65320 39780 65320 39780 0 net158
rlabel metal2 40710 2244 40710 2244 0 net159
rlabel metal1 53406 5134 53406 5134 0 net16
rlabel metal1 63342 45003 63342 45003 0 net160
rlabel metal2 62606 2142 62606 2142 0 net161
rlabel metal2 65412 39644 65412 39644 0 net162
rlabel metal1 29946 2346 29946 2346 0 net163
rlabel metal1 63342 36303 63342 36303 0 net164
rlabel metal1 39284 2618 39284 2618 0 net165
rlabel metal1 63618 45254 63618 45254 0 net166
rlabel metal1 37720 2618 37720 2618 0 net167
rlabel metal1 63342 45731 63342 45731 0 net168
rlabel metal1 32338 2278 32338 2278 0 net169
rlabel metal2 55246 3740 55246 3740 0 net17
rlabel metal1 63986 43826 63986 43826 0 net170
rlabel metal1 67896 1258 67896 1258 0 net171
rlabel metal1 65642 36346 65642 36346 0 net172
rlabel metal1 66056 2618 66056 2618 0 net173
rlabel metal1 63342 72262 63342 72262 0 net174
rlabel metal1 36524 2618 36524 2618 0 net175
rlabel metal1 63618 45948 63618 45948 0 net176
rlabel metal2 32798 3876 32798 3876 0 net177
rlabel metal1 63342 47187 63342 47187 0 net178
rlabel metal1 27094 3536 27094 3536 0 net179
rlabel metal2 55982 3570 55982 3570 0 net18
rlabel metal1 63894 47702 63894 47702 0 net180
rlabel metal1 29532 3162 29532 3162 0 net181
rlabel metal1 63250 47445 63250 47445 0 net182
rlabel metal1 28566 2822 28566 2822 0 net183
rlabel metal2 53774 5015 53774 5015 0 net184
rlabel metal1 28060 3026 28060 3026 0 net185
rlabel metal1 27646 1938 27646 1938 0 net186
rlabel metal1 63342 37517 63342 37517 0 net187
rlabel metal1 26956 2618 26956 2618 0 net188
rlabel metal1 30268 1326 30268 1326 0 net189
rlabel metal1 48714 2516 48714 2516 0 net19
rlabel metal1 63342 55734 63342 55734 0 net190
rlabel metal1 26818 1326 26818 1326 0 net191
rlabel metal1 32752 1326 32752 1326 0 net192
rlabel metal1 63342 82224 63342 82224 0 net193
rlabel metal1 30590 1292 30590 1292 0 net194
rlabel metal2 49450 2244 49450 2244 0 net195
rlabel metal1 49312 1326 49312 1326 0 net196
rlabel metal2 46966 2244 46966 2244 0 net197
rlabel metal1 46414 1394 46414 1394 0 net198
rlabel metal1 45264 2074 45264 2074 0 net199
rlabel metal2 41354 3366 41354 3366 0 net2
rlabel metal1 61502 2040 61502 2040 0 net20
rlabel metal2 43010 2652 43010 2652 0 net200
rlabel metal2 41446 2244 41446 2244 0 net201
rlabel metal1 39928 1870 39928 1870 0 net202
rlabel metal2 37858 2788 37858 2788 0 net203
rlabel metal1 35558 1530 35558 1530 0 net204
rlabel metal1 53912 1326 53912 1326 0 net205
rlabel metal1 32338 2380 32338 2380 0 net206
rlabel metal1 56534 1326 56534 1326 0 net207
rlabel metal2 52670 2244 52670 2244 0 net208
rlabel metal2 55614 2244 55614 2244 0 net209
rlabel metal1 62790 2584 62790 2584 0 net21
rlabel metal2 60030 2108 60030 2108 0 net210
rlabel metal2 50830 1802 50830 1802 0 net211
rlabel metal1 59616 1326 59616 1326 0 net212
rlabel metal1 33396 2414 33396 2414 0 net213
rlabel metal2 61410 2244 61410 2244 0 net214
rlabel metal1 62146 1326 62146 1326 0 net215
rlabel metal1 28060 3162 28060 3162 0 net216
rlabel metal1 30452 2822 30452 2822 0 net217
rlabel metal1 65504 1258 65504 1258 0 net218
rlabel metal1 66516 1870 66516 1870 0 net219
rlabel metal1 64860 1496 64860 1496 0 net22
rlabel metal1 26864 1870 26864 1870 0 net220
rlabel metal1 67436 2958 67436 2958 0 net221
rlabel metal1 65044 2822 65044 2822 0 net222
rlabel metal1 24932 1870 24932 1870 0 net223
rlabel metal1 69552 1530 69552 1530 0 net224
rlabel metal1 69920 2074 69920 2074 0 net225
rlabel metal1 73324 1326 73324 1326 0 net226
rlabel metal1 43884 2414 43884 2414 0 net227
rlabel metal1 43286 1326 43286 1326 0 net228
rlabel metal2 41262 1734 41262 1734 0 net229
rlabel metal1 62077 1734 62077 1734 0 net23
rlabel metal1 38456 1530 38456 1530 0 net230
rlabel metal2 37030 2244 37030 2244 0 net231
rlabel metal1 30958 1530 30958 1530 0 net232
rlabel metal2 36018 2652 36018 2652 0 net233
rlabel metal1 31832 2618 31832 2618 0 net234
rlabel metal1 29716 2618 29716 2618 0 net235
rlabel metal1 26312 2074 26312 2074 0 net236
rlabel via1 33166 2805 33166 2805 0 net24
rlabel metal2 62698 2278 62698 2278 0 net25
rlabel metal1 66608 31790 66608 31790 0 net26
rlabel metal1 66516 32878 66516 32878 0 net27
rlabel metal1 63894 2278 63894 2278 0 net28
rlabel metal1 63618 1768 63618 1768 0 net29
rlabel metal1 55154 3128 55154 3128 0 net3
rlabel metal1 67344 36142 67344 36142 0 net30
rlabel metal1 66654 37774 66654 37774 0 net31
rlabel metal1 67850 2006 67850 2006 0 net32
rlabel metal1 67390 39406 67390 39406 0 net33
rlabel metal1 70610 2006 70610 2006 0 net34
rlabel metal2 47610 4522 47610 4522 0 net35
rlabel metal1 70748 2482 70748 2482 0 net36
rlabel metal1 71024 2346 71024 2346 0 net37
rlabel metal1 39054 2550 39054 2550 0 net38
rlabel metal1 34454 4590 34454 4590 0 net39
rlabel metal2 26910 3519 26910 3519 0 net4
rlabel metal1 45402 4760 45402 4760 0 net40
rlabel metal1 40434 3536 40434 3536 0 net41
rlabel metal2 40894 3910 40894 3910 0 net42
rlabel metal1 51428 5678 51428 5678 0 net43
rlabel metal2 51750 4420 51750 4420 0 net44
rlabel metal1 28474 1836 28474 1836 0 net45
rlabel metal2 33994 2210 33994 2210 0 net46
rlabel metal1 31694 1224 31694 1224 0 net47
rlabel metal3 65527 34748 65527 34748 0 net48
rlabel metal2 25162 1870 25162 1870 0 net49
rlabel metal1 28658 4488 28658 4488 0 net5
rlabel metal2 27094 2278 27094 2278 0 net50
rlabel metal2 25714 1156 25714 1156 0 net51
rlabel metal2 28198 2074 28198 2074 0 net52
rlabel metal2 40066 3264 40066 3264 0 net53
rlabel metal1 43240 1938 43240 1938 0 net54
rlabel metal1 33994 986 33994 986 0 net55
rlabel metal2 47518 1088 47518 1088 0 net56
rlabel metal1 33810 1462 33810 1462 0 net57
rlabel metal2 32430 5321 32430 5321 0 net58
rlabel metal1 49772 2006 49772 2006 0 net59
rlabel metal3 66033 12716 66033 12716 0 net6
rlabel metal1 52486 1326 52486 1326 0 net60
rlabel metal1 53314 1938 53314 1938 0 net61
rlabel metal1 55062 1326 55062 1326 0 net62
rlabel metal1 29302 1360 29302 1360 0 net63
rlabel metal1 54556 1938 54556 1938 0 net64
rlabel metal1 57546 2414 57546 2414 0 net65
rlabel metal2 57638 3706 57638 3706 0 net66
rlabel metal2 63664 1326 63664 1326 0 net67
rlabel metal1 63710 2448 63710 2448 0 net68
rlabel metal3 62468 4148 62468 4148 0 net69
rlabel metal2 36294 3961 36294 3961 0 net7
rlabel metal1 63664 3026 63664 3026 0 net70
rlabel metal1 66010 2414 66010 2414 0 net71
rlabel metal1 69092 1938 69092 1938 0 net72
rlabel metal2 69414 3468 69414 3468 0 net73
rlabel metal1 32476 1938 32476 1938 0 net74
rlabel metal1 70656 1326 70656 1326 0 net75
rlabel metal2 71438 2924 71438 2924 0 net76
rlabel metal1 33488 3910 33488 3910 0 net77
rlabel metal1 34040 1938 34040 1938 0 net78
rlabel metal1 35512 1326 35512 1326 0 net79
rlabel metal1 36202 3604 36202 3604 0 net8
rlabel metal1 35926 1938 35926 1938 0 net80
rlabel metal1 37996 3026 37996 3026 0 net81
rlabel metal2 39790 2244 39790 2244 0 net82
rlabel metal1 40894 4012 40894 4012 0 net83
rlabel metal2 35742 4352 35742 4352 0 net84
rlabel metal2 40158 3451 40158 3451 0 net85
rlabel metal1 35052 4590 35052 4590 0 net86
rlabel metal1 40710 4182 40710 4182 0 net87
rlabel metal1 29900 4658 29900 4658 0 net88
rlabel metal1 40710 4046 40710 4046 0 net89
rlabel metal2 37490 3009 37490 3009 0 net9
rlabel metal1 63487 49657 63487 49657 0 net90
rlabel metal1 63342 43713 63342 43713 0 net91
rlabel metal1 63342 42543 63342 42543 0 net92
rlabel metal1 63342 50114 63342 50114 0 net93
rlabel metal1 63441 52094 63441 52094 0 net94
rlabel metal1 63342 52289 63342 52289 0 net95
rlabel metal1 63487 48715 63487 48715 0 net96
rlabel via3 65757 46988 65757 46988 0 net97
rlabel metal3 66079 46988 66079 46988 0 net98
rlabel metal1 48944 2414 48944 2414 0 net99
rlabel metal2 23138 493 23138 493 0 wb_clk_i
rlabel metal2 23506 1044 23506 1044 0 wb_rst_i
rlabel metal2 23966 1078 23966 1078 0 wbs_ack_o
rlabel metal2 41446 874 41446 874 0 wbs_adr_i[10]
rlabel metal2 42826 1588 42826 1588 0 wbs_adr_i[11]
rlabel metal2 25438 1700 25438 1700 0 wbs_adr_i[2]
rlabel metal2 31326 1520 31326 1520 0 wbs_adr_i[3]
rlabel metal2 33166 1078 33166 1078 0 wbs_adr_i[4]
rlabel metal2 29854 1122 29854 1122 0 wbs_adr_i[5]
rlabel metal1 36248 2958 36248 2958 0 wbs_adr_i[6]
rlabel metal2 37306 1316 37306 1316 0 wbs_adr_i[7]
rlabel metal2 38686 1044 38686 1044 0 wbs_adr_i[8]
rlabel metal2 40066 1044 40066 1044 0 wbs_adr_i[9]
rlabel metal2 24426 823 24426 823 0 wbs_cyc_i
rlabel metal2 26266 1622 26266 1622 0 wbs_dat_i[0]
rlabel metal2 41906 823 41906 823 0 wbs_dat_i[10]
rlabel metal2 43286 1282 43286 1282 0 wbs_dat_i[11]
rlabel metal2 44666 976 44666 976 0 wbs_dat_i[12]
rlabel metal2 46046 1316 46046 1316 0 wbs_dat_i[13]
rlabel metal2 47426 1588 47426 1588 0 wbs_dat_i[14]
rlabel metal2 48806 1316 48806 1316 0 wbs_dat_i[15]
rlabel metal2 50186 1588 50186 1588 0 wbs_dat_i[16]
rlabel metal2 51566 1316 51566 1316 0 wbs_dat_i[17]
rlabel metal2 52946 976 52946 976 0 wbs_dat_i[18]
rlabel metal2 54326 823 54326 823 0 wbs_dat_i[19]
rlabel metal2 28106 2404 28106 2404 0 wbs_dat_i[1]
rlabel metal2 55706 976 55706 976 0 wbs_dat_i[20]
rlabel metal2 57086 1350 57086 1350 0 wbs_dat_i[21]
rlabel metal2 58466 1027 58466 1027 0 wbs_dat_i[22]
rlabel metal2 59846 1316 59846 1316 0 wbs_dat_i[23]
rlabel metal2 61226 1044 61226 1044 0 wbs_dat_i[24]
rlabel metal2 62606 1044 62606 1044 0 wbs_dat_i[25]
rlabel metal2 63986 1860 63986 1860 0 wbs_dat_i[26]
rlabel metal2 65366 1316 65366 1316 0 wbs_dat_i[27]
rlabel metal2 66746 1044 66746 1044 0 wbs_dat_i[28]
rlabel metal2 68126 1044 68126 1044 0 wbs_dat_i[29]
rlabel metal1 29348 3026 29348 3026 0 wbs_dat_i[2]
rlabel metal2 69506 874 69506 874 0 wbs_dat_i[30]
rlabel metal2 70886 1044 70886 1044 0 wbs_dat_i[31]
rlabel metal2 31786 1860 31786 1860 0 wbs_dat_i[3]
rlabel metal2 33626 1622 33626 1622 0 wbs_dat_i[4]
rlabel metal2 35006 1588 35006 1588 0 wbs_dat_i[5]
rlabel metal2 36386 1044 36386 1044 0 wbs_dat_i[6]
rlabel metal2 37766 1588 37766 1588 0 wbs_dat_i[7]
rlabel metal2 39146 1316 39146 1316 0 wbs_dat_i[8]
rlabel metal2 40526 1078 40526 1078 0 wbs_dat_i[9]
rlabel metal2 26726 959 26726 959 0 wbs_dat_o[0]
rlabel metal2 42366 891 42366 891 0 wbs_dat_o[10]
rlabel metal2 43746 1316 43746 1316 0 wbs_dat_o[11]
rlabel metal2 45126 1010 45126 1010 0 wbs_dat_o[12]
rlabel metal2 46506 1010 46506 1010 0 wbs_dat_o[13]
rlabel metal2 47886 1316 47886 1316 0 wbs_dat_o[14]
rlabel metal2 49266 1078 49266 1078 0 wbs_dat_o[15]
rlabel metal2 50646 1316 50646 1316 0 wbs_dat_o[16]
rlabel metal2 52026 823 52026 823 0 wbs_dat_o[17]
rlabel metal2 53406 1316 53406 1316 0 wbs_dat_o[18]
rlabel metal2 54786 1010 54786 1010 0 wbs_dat_o[19]
rlabel metal2 28566 1010 28566 1010 0 wbs_dat_o[1]
rlabel metal2 56166 1316 56166 1316 0 wbs_dat_o[20]
rlabel metal2 57546 1622 57546 1622 0 wbs_dat_o[21]
rlabel metal1 58880 3434 58880 3434 0 wbs_dat_o[22]
rlabel metal2 64630 1122 64630 1122 0 wbs_dat_o[23]
rlabel metal2 61686 1520 61686 1520 0 wbs_dat_o[24]
rlabel metal2 63066 891 63066 891 0 wbs_dat_o[25]
rlabel metal2 64446 823 64446 823 0 wbs_dat_o[26]
rlabel metal2 65826 1622 65826 1622 0 wbs_dat_o[27]
rlabel metal2 67206 1316 67206 1316 0 wbs_dat_o[28]
rlabel metal1 69230 2958 69230 2958 0 wbs_dat_o[29]
rlabel metal2 30406 1316 30406 1316 0 wbs_dat_o[2]
rlabel metal2 69966 1078 69966 1078 0 wbs_dat_o[30]
rlabel metal2 71346 1316 71346 1316 0 wbs_dat_o[31]
rlabel metal2 32246 1316 32246 1316 0 wbs_dat_o[3]
rlabel metal2 34086 1316 34086 1316 0 wbs_dat_o[4]
rlabel metal2 35466 823 35466 823 0 wbs_dat_o[5]
rlabel metal2 36846 1282 36846 1282 0 wbs_dat_o[6]
rlabel metal2 38226 823 38226 823 0 wbs_dat_o[7]
rlabel metal2 39606 1010 39606 1010 0 wbs_dat_o[8]
rlabel metal2 40986 1010 40986 1010 0 wbs_dat_o[9]
rlabel metal2 27186 1588 27186 1588 0 wbs_sel_i[0]
rlabel metal1 29118 4046 29118 4046 0 wbs_sel_i[1]
rlabel metal1 26174 1292 26174 1292 0 wbs_sel_i[2]
rlabel metal2 27278 1088 27278 1088 0 wbs_sel_i[3]
rlabel metal2 24886 1588 24886 1588 0 wbs_stb_i
rlabel metal2 25346 1350 25346 1350 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 76000 87000
<< end >>
