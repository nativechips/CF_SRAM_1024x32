magic
tech sky130A
magscale 1 2
timestamp 1578962917
<< checkpaint >>
rect -1260 -1260 78834 62615
<< metal1 >>
rect 38761 61347 38813 61355
rect 38761 61263 38813 61295
rect 1319 0 1365 600
rect 2295 0 2341 600
rect 2547 0 2593 600
rect 3499 0 3545 600
rect 4475 0 4521 600
rect 4727 0 4773 600
rect 5679 0 5725 600
rect 6655 0 6701 600
rect 6907 0 6953 600
rect 7859 0 7905 600
rect 8835 0 8881 600
rect 9087 0 9133 600
rect 10039 0 10085 600
rect 11015 0 11061 600
rect 11267 0 11313 600
rect 12219 0 12265 600
rect 13195 0 13241 600
rect 13447 0 13493 600
rect 14399 0 14445 600
rect 15375 0 15421 600
rect 15627 0 15673 600
rect 16579 0 16625 600
rect 17555 0 17601 600
rect 17807 0 17853 600
rect 18759 0 18805 600
rect 19735 0 19781 600
rect 19987 0 20033 600
rect 20939 0 20985 600
rect 21915 0 21961 600
rect 22167 0 22213 600
rect 23119 0 23165 600
rect 24095 0 24141 600
rect 24347 0 24393 600
rect 25299 0 25345 600
rect 26275 0 26321 600
rect 26527 0 26573 600
rect 27479 0 27525 600
rect 28455 0 28501 600
rect 28707 0 28753 600
rect 29659 0 29705 600
rect 30635 0 30681 600
rect 30887 0 30933 600
rect 31839 0 31885 600
rect 32815 0 32861 600
rect 33067 0 33113 600
rect 34019 0 34065 600
rect 34383 0 34421 600
rect 34995 0 35041 600
rect 35247 0 35293 600
rect 35628 0 35680 600
rect 35813 0 35865 600
rect 36441 0 36493 600
rect 36521 0 36573 600
rect 37149 0 37201 601
rect 37229 0 37281 600
rect 37857 0 37909 601
rect 37937 0 37989 600
rect 39273 0 39325 600
rect 39353 0 39405 600
rect 39981 0 40033 600
rect 40061 0 40113 600
rect 40689 496 40741 735
rect 40689 0 40741 444
rect 40769 0 40821 600
rect 41637 0 41677 600
rect 41705 0 41745 600
rect 41977 0 42015 600
rect 42281 0 42327 600
rect 42533 0 42579 600
rect 43509 0 43555 600
rect 44069 0 44119 600
rect 44147 0 44195 600
rect 44461 0 44507 600
rect 44713 0 44759 600
rect 45409 0 45455 600
rect 45689 0 45735 600
rect 46641 0 46687 600
rect 46893 0 46939 600
rect 47869 0 47915 600
rect 48821 0 48867 600
rect 49073 0 49119 600
rect 50049 0 50095 600
rect 51001 0 51047 600
rect 51253 0 51299 600
rect 52229 0 52275 600
rect 53181 0 53227 600
rect 53433 0 53479 600
rect 54409 0 54455 600
rect 55361 0 55407 600
rect 55613 0 55659 600
rect 56589 0 56635 600
rect 57541 0 57587 600
rect 57793 0 57839 600
rect 58769 0 58815 600
rect 59721 0 59767 600
rect 59973 0 60019 600
rect 60949 0 60995 600
rect 61901 0 61947 600
rect 62153 0 62199 600
rect 63129 0 63175 600
rect 64081 0 64127 600
rect 64333 0 64379 600
rect 65309 0 65355 600
rect 66261 0 66307 600
rect 66513 0 66559 600
rect 67489 0 67535 600
rect 68441 0 68487 600
rect 68693 0 68739 600
rect 69669 0 69715 600
rect 70621 0 70667 600
rect 70873 0 70919 600
rect 71849 0 71895 600
rect 72801 0 72847 600
rect 73053 0 73099 600
rect 74029 0 74075 600
rect 74981 0 75027 600
rect 75233 0 75279 600
rect 76209 0 76255 600
<< via1 >>
rect 38761 61295 38813 61347
rect 40689 444 40741 496
<< metal2 >>
rect 38750 61293 38759 61349
rect 38815 61293 38824 61349
rect 0 60810 56 61263
rect 228 61159 77346 61263
rect 356 60931 77218 61131
rect 77518 60810 77574 61263
rect 602 57815 76972 57909
rect 246 57668 77328 57762
rect 602 54925 76972 55019
rect 246 54778 77328 54872
rect 602 52035 76972 52129
rect 246 51888 77328 51982
rect 602 49145 76972 49239
rect 246 48998 77328 49092
rect 602 46255 76972 46349
rect 246 46108 77328 46202
rect 602 43365 76972 43459
rect 246 43218 77328 43312
rect 602 40475 76972 40569
rect 246 40328 77328 40422
rect 602 37585 76972 37679
rect 246 37438 77328 37532
rect 602 34695 76972 34789
rect 246 34548 77328 34642
rect 602 31805 76972 31899
rect 246 31658 77328 31752
rect 602 28915 76972 29009
rect 246 28768 77328 28862
rect 602 26025 76972 26119
rect 246 25878 77328 25972
rect 602 23135 76972 23229
rect 246 22988 77328 23082
rect 602 20245 76972 20339
rect 246 20098 77328 20192
rect 602 17355 76972 17449
rect 246 17208 77328 17302
rect 356 14408 35816 14502
rect 41758 14408 77218 14502
rect 228 14200 35816 14294
rect 41758 14200 77346 14294
rect 196 13453 35816 13653
rect 41758 13453 77378 13653
rect 0 11572 196 13241
rect 77378 11572 77574 13241
rect 806 10963 76768 11073
rect 0 10452 192 10888
rect 77382 10452 77574 10888
rect 806 10235 35686 10363
rect 41888 10235 76768 10363
rect 780 10077 76794 10205
rect 0 9013 192 9768
rect 806 9721 76768 9849
rect 806 9553 76768 9681
rect 806 9385 35686 9513
rect 41888 9385 76768 9513
rect 77382 9013 77574 9768
rect 806 8641 76768 8769
rect 806 8403 76768 8531
rect 0 7907 192 8329
rect 806 8257 76768 8373
rect 806 7810 76768 7938
rect 77382 7907 77574 8329
rect 806 7535 76768 7663
rect 0 6862 192 7223
rect 806 6957 76768 7085
rect 77382 6862 77574 7223
rect 806 6664 76768 6792
rect 806 6518 76768 6634
rect 806 6214 76768 6330
rect 0 5862 192 6178
rect 77382 5862 77574 6178
rect 806 5372 76768 5488
rect 0 4862 192 5178
rect 806 5162 76768 5342
rect 35686 4874 41888 4938
rect 806 4822 76768 4874
rect 77382 4862 77574 5178
rect 806 4758 35686 4822
rect 41888 4758 76768 4822
rect 806 4149 76768 4265
rect 0 4047 192 4099
rect 806 3979 76768 4119
rect 77382 4047 77574 4099
rect 806 3833 76768 3949
rect 0 3671 192 3723
rect 77382 3671 77574 3723
rect 806 3525 76768 3641
rect 806 3379 76768 3495
rect 806 3173 76768 3349
rect 806 3149 35686 3173
rect 41888 3149 76768 3173
rect 0 2671 192 2987
rect 806 2871 76768 2987
rect 806 2859 35686 2871
rect 41888 2859 76768 2871
rect 806 2713 76768 2829
rect 77382 2671 77574 2987
rect 0 1671 192 1987
rect 77382 1671 77574 1987
rect 0 672 192 987
rect 806 802 76768 976
rect 806 600 76768 774
rect 77382 672 77574 987
rect 38750 442 38759 498
rect 38815 484 38824 498
rect 40683 484 40689 496
rect 38815 456 40689 484
rect 38815 442 38824 456
rect 40683 444 40689 456
rect 40741 444 40747 496
<< via2 >>
rect 38759 61347 38815 61349
rect 38759 61295 38761 61347
rect 38761 61295 38813 61347
rect 38813 61295 38815 61347
rect 38759 61293 38815 61295
rect 38759 442 38815 498
<< metal3 >>
rect 38754 61349 38820 61354
rect 38754 61293 38759 61349
rect 38815 61293 38820 61349
rect 38754 61288 38820 61293
rect 38757 503 38817 61288
rect 38754 498 38820 503
rect 38754 442 38759 498
rect 38815 442 38820 498
rect 38754 437 38820 442
use CF_SRAM_1024x32  CF_SRAM_1024x32_macro_0
timestamp 1578962917
transform 1 0 0 0 1 600
box 0 0 77574 60663
<< labels >>
rlabel metal1 s 40689 600 40741 735 4 WLOFF
port 2 nsew
rlabel metal1 s 40715 667 40715 667 4 WLOFF
rlabel metal1 s 40689 0 40741 400 4 WLOFF
port 2 nsew
rlabel metal1 s 42281 0 42327 400 4 DO[16]
port 3 nsew
rlabel metal1 s 43509 0 43555 400 4 BEN[16]
port 4 nsew
rlabel metal1 s 44461 0 44507 400 4 DO[17]
port 5 nsew
rlabel metal1 s 45689 0 45735 400 4 BEN[17]
port 6 nsew
rlabel metal1 s 46641 0 46687 400 4 DO[18]
port 7 nsew
rlabel metal1 s 47869 0 47915 400 4 BEN[18]
port 8 nsew
rlabel metal1 s 48821 0 48867 400 4 DO[19]
port 9 nsew
rlabel metal1 s 50049 0 50095 400 4 BEN[19]
port 10 nsew
rlabel metal1 s 51001 0 51047 400 4 DO[20]
port 11 nsew
rlabel metal1 s 52229 0 52275 400 4 BEN[20]
port 12 nsew
rlabel metal1 s 53181 0 53227 400 4 DO[21]
port 13 nsew
rlabel metal1 s 54409 0 54455 400 4 BEN[21]
port 14 nsew
rlabel metal1 s 55361 0 55407 400 4 DO[22]
port 15 nsew
rlabel metal1 s 56589 0 56635 400 4 BEN[22]
port 16 nsew
rlabel metal1 s 57541 0 57587 400 4 DO[23]
port 17 nsew
rlabel metal1 s 58769 0 58815 400 4 BEN[23]
port 18 nsew
rlabel metal1 s 59721 0 59767 400 4 DO[24]
port 19 nsew
rlabel metal1 s 60949 0 60995 400 4 BEN[24]
port 20 nsew
rlabel metal1 s 61901 0 61947 400 4 DO[25]
port 21 nsew
rlabel metal1 s 63129 0 63175 400 4 BEN[25]
port 22 nsew
rlabel metal1 s 64081 0 64127 400 4 DO[26]
port 23 nsew
rlabel metal1 s 65309 0 65355 400 4 BEN[26]
port 24 nsew
rlabel metal1 s 66261 0 66307 400 4 DO[27]
port 25 nsew
rlabel metal1 s 67489 0 67535 400 4 BEN[27]
port 26 nsew
rlabel metal1 s 68441 0 68487 400 4 DO[28]
port 27 nsew
rlabel metal1 s 69669 0 69715 400 4 BEN[28]
port 28 nsew
rlabel metal1 s 70621 0 70667 400 4 DO[29]
port 29 nsew
rlabel metal1 s 71849 0 71895 400 4 BEN[29]
port 30 nsew
rlabel metal1 s 72801 0 72847 400 4 DO[30]
port 31 nsew
rlabel metal1 s 74029 0 74075 400 4 BEN[30]
port 32 nsew
rlabel metal1 s 74981 0 75027 400 4 DO[31]
port 33 nsew
rlabel metal1 s 76209 0 76255 400 4 BEN[31]
port 34 nsew
rlabel metal1 s 39981 0 40033 400 4 AD[0]
port 35 nsew
rlabel metal1 s 39353 0 39405 400 4 AD[1]
port 36 nsew
rlabel metal1 s 39273 0 39325 400 4 AD[2]
port 37 nsew
rlabel metal1 s 44147 0 44195 400 4 WLBI
port 38 nsew
rlabel metal1 s 45409 0 45455 400 4 CLKin
port 39 nsew
rlabel metal1 s 40769 0 40821 400 4 EN
port 40 nsew
rlabel metal1 s 40061 0 40113 400 4 R_WB
port 41 nsew
rlabel metal1 s 41637 0 41677 400 4 SM
port 42 nsew
rlabel metal1 s 44069 0 44119 400 4 TM
port 43 nsew
rlabel metal1 s 41977 0 42015 400 4 ScanInDR
port 44 nsew
rlabel metal1 s 41705 0 41745 400 4 ScanOutCC
port 45 nsew
rlabel metal1 s 34383 0 34421 400 4 ScanInDL
port 46 nsew
rlabel metal1 s 15627 0 15673 400 4 DO[9]
port 47 nsew
rlabel metal1 s 14399 0 14445 400 4 BEN[9]
port 48 nsew
rlabel metal1 s 13447 0 13493 400 4 DO[10]
port 49 nsew
rlabel metal1 s 12219 0 12265 400 4 BEN[10]
port 50 nsew
rlabel metal1 s 11267 0 11313 400 4 DO[11]
port 51 nsew
rlabel metal1 s 10039 0 10085 400 4 BEN[11]
port 52 nsew
rlabel metal1 s 9087 0 9133 400 4 DO[12]
port 53 nsew
rlabel metal1 s 7859 0 7905 400 4 BEN[12]
port 54 nsew
rlabel metal1 s 6907 0 6953 400 4 DO[13]
port 55 nsew
rlabel metal1 s 5679 0 5725 400 4 BEN[13]
port 56 nsew
rlabel metal1 s 4727 0 4773 400 4 DO[14]
port 57 nsew
rlabel metal1 s 3499 0 3545 400 4 BEN[14]
port 58 nsew
rlabel metal1 s 2547 0 2593 400 4 DO[15]
port 59 nsew
rlabel metal1 s 1319 0 1365 400 4 BEN[15]
port 60 nsew
rlabel metal1 s 16579 0 16625 400 4 BEN[8]
port 61 nsew
rlabel metal1 s 35813 0 35865 400 4 AD[3]
port 62 nsew
rlabel metal1 s 37937 0 37989 400 4 AD[4]
port 63 nsew
rlabel metal1 s 37857 1 37909 400 4 AD[5]
port 64 nsew
rlabel metal1 s 37229 0 37281 400 4 AD[6]
port 65 nsew
rlabel metal1 s 37149 1 37201 400 4 AD[7]
port 66 nsew
rlabel metal1 s 36521 0 36573 400 4 AD[8]
port 67 nsew
rlabel metal1 s 36441 0 36493 400 4 AD[9]
port 68 nsew
rlabel metal1 s 35628 0 35680 400 4 ScanInCC
port 69 nsew
rlabel metal1 s 35247 0 35293 400 4 DO[0]
port 70 nsew
rlabel metal1 s 34019 0 34065 400 4 BEN[0]
port 71 nsew
rlabel metal1 s 33067 0 33113 400 4 DO[1]
port 72 nsew
rlabel metal1 s 31839 0 31885 400 4 BEN[1]
port 73 nsew
rlabel metal1 s 30887 0 30933 400 4 DO[2]
port 74 nsew
rlabel metal1 s 29659 0 29705 400 4 BEN[2]
port 75 nsew
rlabel metal1 s 28707 0 28753 400 4 DO[3]
port 76 nsew
rlabel metal1 s 27479 0 27525 400 4 BEN[3]
port 77 nsew
rlabel metal1 s 26527 0 26573 400 4 DO[4]
port 78 nsew
rlabel metal1 s 25299 0 25345 400 4 BEN[4]
port 79 nsew
rlabel metal1 s 24347 0 24393 400 4 DO[5]
port 80 nsew
rlabel metal1 s 23119 0 23165 400 4 BEN[5]
port 81 nsew
rlabel metal1 s 22167 0 22213 400 4 DO[6]
port 82 nsew
rlabel metal1 s 20939 0 20985 400 4 BEN[6]
port 83 nsew
rlabel metal1 s 19987 0 20033 400 4 DO[7]
port 84 nsew
rlabel metal1 s 18759 0 18805 400 4 BEN[7]
port 85 nsew
rlabel metal1 s 17807 0 17853 400 4 DO[8]
port 86 nsew
rlabel metal1 s 28455 0 28501 400 4 DI[3]
port 87 nsew
rlabel metal1 s 8835 0 8881 400 4 DI[12]
port 88 nsew
rlabel metal1 s 34995 0 35041 400 4 DI[0]
port 89 nsew
rlabel metal1 s 26275 0 26321 400 4 DI[4]
port 90 nsew
rlabel metal1 s 4475 0 4521 400 4 DI[14]
port 91 nsew
rlabel metal1 s 11015 0 11061 400 4 DI[11]
port 92 nsew
rlabel metal1 s 24095 0 24141 400 4 DI[5]
port 93 nsew
rlabel metal1 s 32815 0 32861 400 4 DI[1]
port 94 nsew
rlabel metal1 s 15375 0 15421 400 4 DI[9]
port 95 nsew
rlabel metal1 s 21915 0 21961 400 4 DI[6]
port 96 nsew
rlabel metal1 s 2295 0 2341 400 4 DI[15]
port 97 nsew
rlabel metal1 s 30635 0 30681 400 4 DI[2]
port 98 nsew
rlabel metal1 s 19735 0 19781 400 4 DI[7]
port 99 nsew
rlabel metal1 s 6655 0 6701 400 4 DI[13]
port 100 nsew
rlabel metal1 s 13195 0 13241 400 4 DI[10]
port 101 nsew
rlabel metal1 s 17555 0 17601 400 4 DI[8]
port 102 nsew
rlabel metal1 s 57793 0 57839 400 4 DI[23]
port 103 nsew
rlabel metal1 s 66513 0 66559 400 4 DI[27]
port 104 nsew
rlabel metal1 s 49073 0 49119 400 4 DI[19]
port 105 nsew
rlabel metal1 s 53433 0 53479 400 4 DI[21]
port 106 nsew
rlabel metal1 s 68693 0 68739 400 4 DI[28]
port 107 nsew
rlabel metal1 s 59973 0 60019 400 4 DI[24]
port 108 nsew
rlabel metal1 s 46893 0 46939 400 4 DI[18]
port 109 nsew
rlabel metal1 s 70873 0 70919 400 4 DI[29]
port 110 nsew
rlabel metal1 s 42533 0 42579 400 4 DI[16]
port 111 nsew
rlabel metal1 s 62153 0 62199 400 4 DI[25]
port 112 nsew
rlabel metal1 s 73053 0 73099 400 4 DI[30]
port 113 nsew
rlabel metal1 s 55613 0 55659 400 4 DI[22]
port 114 nsew
rlabel metal1 s 51253 0 51299 400 4 DI[20]
port 115 nsew
rlabel metal1 s 64333 0 64379 400 4 DI[26]
port 116 nsew
rlabel metal1 s 44713 0 44759 400 4 DI[17]
port 117 nsew
rlabel metal1 s 75233 0 75279 400 4 DI[31]
port 118 nsew
rlabel metal2 s 77518 60810 77574 61263 4 vgnd
port 123 nsew
rlabel metal2 s 246 54778 77328 54872 4 vnb
port 119 nsew
rlabel metal2 s 246 51888 77328 51982 4 vnb
port 119 nsew
rlabel metal2 s 246 48998 77328 49092 4 vnb
port 119 nsew
rlabel metal2 s 246 46108 77328 46202 4 vnb
port 119 nsew
rlabel metal2 s 246 43218 77328 43312 4 vnb
port 119 nsew
rlabel metal2 s 246 40328 77328 40422 4 vnb
port 119 nsew
rlabel metal2 s 246 37438 77328 37532 4 vnb
port 119 nsew
rlabel metal2 s 246 34548 77328 34642 4 vnb
port 119 nsew
rlabel metal2 s 246 31658 77328 31752 4 vnb
port 119 nsew
rlabel metal2 s 356 60931 77218 61131 4 vpwra
port 121 nsew
rlabel metal2 s 228 61159 77346 61263 4 vgnd
port 123 nsew
rlabel metal2 s 246 57668 77328 57762 4 vnb
port 119 nsew
rlabel metal2 s 0 60810 56 61263 4 vgnd
port 123 nsew
rlabel metal2 s 602 57815 76972 57909 4 vpb
port 124 nsew
rlabel metal2 s 602 54925 76972 55019 4 vpb
port 124 nsew
rlabel metal2 s 602 52035 76972 52129 4 vpb
port 124 nsew
rlabel metal2 s 602 49145 76972 49239 4 vpb
port 124 nsew
rlabel metal2 s 602 46255 76972 46349 4 vpb
port 124 nsew
rlabel metal2 s 602 43365 76972 43459 4 vpb
port 124 nsew
rlabel metal2 s 602 40475 76972 40569 4 vpb
port 124 nsew
rlabel metal2 s 602 37585 76972 37679 4 vpb
port 124 nsew
rlabel metal2 s 602 34695 76972 34789 4 vpb
port 124 nsew
rlabel metal2 s 602 31805 76972 31899 4 vpb
port 124 nsew
rlabel metal2 s 356 14408 35816 14502 4 vpwra
port 121 nsew
rlabel metal2 s 0 10452 192 10888 4 vpwra
port 121 nsew
rlabel metal2 s 806 3979 76768 4119 4 vpwra
port 121 nsew
rlabel metal2 s 196 13453 35816 13653 4 vpwrp
port 122 nsew
rlabel metal2 s 0 11572 196 13241 4 vpwrp
port 122 nsew
rlabel metal2 s 806 10235 35686 10363 4 vpwrp
port 122 nsew
rlabel metal2 s 806 9721 76768 9849 4 vpwrp
port 122 nsew
rlabel metal2 s 806 8403 76768 8531 4 vpwrp
port 122 nsew
rlabel metal2 s 0 7907 192 8329 4 vpwrp
port 122 nsew
rlabel metal2 s 806 7810 76768 7938 4 vpwrp
port 122 nsew
rlabel metal2 s 806 6664 76768 6792 4 vpwrp
port 122 nsew
rlabel metal2 s 806 5162 76768 5342 4 vpwrp
port 122 nsew
rlabel metal2 s 0 4862 192 5178 4 vpwrp
port 122 nsew
rlabel metal2 s 806 3833 76768 3949 4 vpwrp
port 122 nsew
rlabel metal2 s 806 3379 76768 3495 4 vpwrp
port 122 nsew
rlabel metal2 s 806 802 76768 976 4 vpwrp
port 122 nsew
rlabel metal2 s 0 672 192 987 4 vpwrp
port 122 nsew
rlabel metal2 s 0 4047 192 4099 4 vpwrac
port 126 nsew
rlabel metal2 s 246 28768 77328 28862 4 vnb
port 119 nsew
rlabel metal2 s 246 25878 77328 25972 4 vnb
port 119 nsew
rlabel metal2 s 228 14200 35816 14294 4 vgnd
port 123 nsew
rlabel metal2 s 806 10963 76768 11073 4 vgnd
port 123 nsew
rlabel metal2 s 806 9553 76768 9681 4 vgnd
port 123 nsew
rlabel metal2 s 0 9013 192 9768 4 vgnd
port 123 nsew
rlabel metal2 s 806 8641 76768 8769 4 vgnd
port 123 nsew
rlabel metal2 s 806 8257 76768 8373 4 vgnd
port 123 nsew
rlabel metal2 s 806 7535 76768 7663 4 vgnd
port 123 nsew
rlabel metal2 s 806 6957 76768 7085 4 vgnd
port 123 nsew
rlabel metal2 s 806 6518 76768 6634 4 vgnd
port 123 nsew
rlabel metal2 s 806 6214 76768 6330 4 vgnd
port 123 nsew
rlabel metal2 s 0 5862 192 6178 4 vgnd
port 123 nsew
rlabel metal2 s 806 5372 76768 5488 4 vgnd
port 123 nsew
rlabel metal2 s 806 4822 76768 4874 4 vgnd
port 123 nsew
rlabel metal2 s 806 4758 35686 4822 4 vgnd
port 123 nsew
rlabel metal2 s 35686 4874 41888 4938 4 vgnd
port 123 nsew
rlabel metal2 s 806 4149 76768 4265 4 vgnd
port 123 nsew
rlabel metal2 s 806 2713 76768 2829 4 vgnd
port 123 nsew
rlabel metal2 s 0 1671 192 1987 4 vgnd
port 123 nsew
rlabel metal2 s 806 600 76768 774 4 vgnd
port 123 nsew
rlabel metal2 s 246 22988 77328 23082 4 vnb
port 119 nsew
rlabel metal2 s 246 20098 77328 20192 4 vnb
port 119 nsew
rlabel metal2 s 246 17208 77328 17302 4 vnb
port 119 nsew
rlabel metal2 s 806 9385 35686 9513 4 vnb
port 119 nsew
rlabel metal2 s 806 2871 76768 2987 4 vnb
port 119 nsew
rlabel metal2 s 806 2859 35686 2871 4 vnb
port 119 nsew
rlabel metal2 s 0 2671 192 2987 4 vnb
port 119 nsew
rlabel metal2 s 806 3173 76768 3349 4 vpwrm
port 120 nsew
rlabel metal2 s 806 3149 35686 3173 4 vpwrm
port 120 nsew
rlabel metal2 s 0 3671 192 3723 4 vpwrpc
port 125 nsew
rlabel metal2 s 602 28915 76972 29009 4 vpb
port 124 nsew
rlabel metal2 s 602 26025 76972 26119 4 vpb
port 124 nsew
rlabel metal2 s 602 23135 76972 23229 4 vpb
port 124 nsew
rlabel metal2 s 602 20245 76972 20339 4 vpb
port 124 nsew
rlabel metal2 s 602 17355 76972 17449 4 vpb
port 124 nsew
rlabel metal2 s 780 10077 76794 10205 4 vpb
port 124 nsew
rlabel metal2 s 0 6862 192 7223 4 vpb
port 124 nsew
rlabel metal2 s 806 3525 76768 3641 4 vpb
port 124 nsew
rlabel metal2 s 77382 9013 77574 9768 4 vgnd
port 123 nsew
rlabel metal2 s 41758 13453 77378 13653 4 vpwrp
port 122 nsew
rlabel metal2 s 77382 4862 77574 5178 4 vpwrp
port 122 nsew
rlabel metal2 s 41888 2859 76768 2871 4 vnb
port 119 nsew
rlabel metal2 s 41888 3149 76768 3173 4 vpwrm
port 120 nsew
rlabel metal2 s 77378 11572 77574 13241 4 vpwrp
port 122 nsew
rlabel metal2 s 77382 3671 77574 3723 4 vpwrpc
port 125 nsew
rlabel metal2 s 41888 10235 76768 10363 4 vpwrp
port 122 nsew
rlabel metal2 s 77382 672 77574 987 4 vpwrp
port 122 nsew
rlabel metal2 s 77382 5862 77574 6178 4 vgnd
port 123 nsew
rlabel metal2 s 77382 2671 77574 2987 4 vnb
port 119 nsew
rlabel metal2 s 41758 14408 77218 14502 4 vpwra
port 121 nsew
rlabel metal2 s 41888 4758 76768 4822 4 vgnd
port 123 nsew
rlabel metal2 s 77382 7907 77574 8329 4 vpwrp
port 122 nsew
rlabel metal2 s 41758 14200 77346 14294 4 vgnd
port 123 nsew
rlabel metal2 s 41888 9385 76768 9513 4 vnb
port 119 nsew
rlabel metal2 s 77382 10452 77574 10888 4 vpwra
port 121 nsew
rlabel metal2 s 77382 6862 77574 7223 4 vpb
port 124 nsew
rlabel metal2 s 77382 4047 77574 4099 4 vpwrac
port 126 nsew
rlabel metal2 s 77382 1671 77574 1987 4 vgnd
port 123 nsew
<< properties >>
string FIXED_BBOX 0 0 77574 61355
<< end >>
